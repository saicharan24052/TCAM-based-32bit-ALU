`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/05/2024 11:28:18 AM
// Design Name: 
// Module Name: multiplier_un
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adder_4bit_re(
input bit clk,
  input logic write_en,
  input logic [3:0] a, b, c,
  input logic [2:0] data_add [63:0],
  input logic [4:0] data_unq [127:0],
  output logic [5:0] sum, actual_sum,
  output logic [12:0] address

    );
    
 logic [4:0] cam_mem [127:0]; // CAM cell 
  logic [2:0] cam_mem_add [63:0]; // CAM cell 
      logic match_flag_0, match_flag_1, match_flag_2, match_flag_3,match_flag_4;
      logic match_flag_carry_1, match_flag_carry_2, match_flag_carry_3,match_flag_carry_4;
      logic data_flag,data_flag_1, sum_flag; 
      int i,i1, j, k, l, m, n, o, p, q, r;
      int addr_0, addr_1, addr_2, addr_3, pp1;
      logic [5:0] sum_reg;
      logic [5:0] late_0,late_1,late_2;
      
      
      /////////   writing data into cam_mem ///////////////////////
       always_ff @(posedge clk) begin 
         if (write_en) begin
           for (i = 0; i < 128; i++) begin
             cam_mem[i] = data_unq[i];
            
           end
           data_flag = 1'b1;
         end 
       end
       
             always_ff @(posedge clk) begin 
         if (write_en) begin
           for (i1 = 0; i1 < 8; i1++) begin
             cam_mem_add[i1] = data_add[i1];
            
           end
           data_flag_1 = 1'b1;
         end 
       end 
       
     //////  end    //////////////////////////////////  
     
     
     
 ///////////////  stage 1   /////////////////////    
     always_ff @(posedge clk) begin 
         if (data_flag) begin 
           match_flag_0 = 1'b0;
           addr_0 = 3'b0;
           
           for (j = 0; j < 8; j++ ) begin  
             if ({a[0], b[0], c[0]} == j[2:0]) begin
               match_flag_0 = 1'b1;
               addr_0 = j[2:0];
               break; // exit the loop once a match is found
             end
           end
         end 
       end       
         
       always_ff @(posedge clk) begin 
         if (data_flag) begin 
           match_flag_1 = 1'b0;
           addr_1 = 3'b0;
           
           for (k = 0; k < 8; k++ ) begin  
             if ({a[1], b[1], c[1]} == k[2:0]) begin
               match_flag_1 = 1'b1;
               addr_1 = k[2:0];
               break; // exit the loop once a match is found
             end
           end
         end 
       end       
     
       always_ff @(posedge clk) begin 
         if (data_flag) begin 
           match_flag_2 = 1'b0;
           addr_2 = 3'b0;
           
           for (l = 0; l < 8; l++ ) begin  
             if ({a[2], b[2], c[2]} == l[2:0]) begin
               match_flag_2 = 1'b1;
               addr_2 = l[2:0];
               break; // exit the loop once a match is found
             end
           end
         end 
       end   
       
       always_ff @(posedge clk) begin 
         if (data_flag) begin 
           match_flag_3 = 1'b0;
           addr_3 = 3'b0;
           
           for (m = 0; m < 8; m++ ) begin  
             if ({a[3], b[3], c[3]} == m[2:0]) begin
               match_flag_3 = 1'b1;
               addr_3 = m[2:0];
               break; // exit the loop once a match is found
             end
           end
         end 
       end   
       
  ///////////////  end  of  stage 1   /////////////////////          
  
  
  always_comb begin
    sum_flag = 1'b0;
    if (match_flag_0 && match_flag_1 && match_flag_2 && match_flag_3) begin
      sum_flag = 1'b1;
    end
  end
  
  
  ///////////////  stage 2   /////////////////////        
  
    always_ff @(posedge clk) begin 
    if (sum_flag) begin 
      match_flag_carry_1 = 1'b0;
      match_flag_carry_2 = 1'b0;
      match_flag_carry_3 = 1'b0;
      match_flag_carry_4 = 1'b0;
      pp1 = 3'b0;
      
     if( {cam_mem_add[addr_3][0], cam_mem_add[addr_2][0]} == 2'b00) begin
          for (n = 0; n < 32; n = n + 1) begin  
              if ({cam_mem_add[addr_1][0], cam_mem_add[addr_3][1], cam_mem_add[addr_2][1], cam_mem_add[addr_1][1], cam_mem_add[addr_0][1]} ==  n[4:0]) begin
                  match_flag_carry_1 = 1'b1;
                  pp1 = {2'b00, n[4:0]};
                  break; // exit the loop once a match is found
              end
          end
      end
      
      if( {cam_mem_add[addr_3][0], cam_mem_add[addr_2][0]} == 2'b01) begin
          for (o = 0; o < 32; o = o + 1) begin  
              if ({cam_mem_add[addr_1][0], cam_mem_add[addr_3][1], cam_mem_add[addr_2][1], cam_mem_add[addr_1][1], cam_mem_add[addr_0][1]} ==  o[4:0]) begin
                  match_flag_carry_2 = 1'b1;
                  pp1 = {2'b01, o[4:0]};
                  break; // exit the loop once a match is found
              end
          end
      end
      
      if( {cam_mem_add[addr_3][0], cam_mem_add[addr_2][0]} == 2'b10) begin
          for (p = 0; p < 32; p = p + 1) begin  
              if ({cam_mem_add[addr_1][0], cam_mem_add[addr_3][1], cam_mem_add[addr_2][1], cam_mem_add[addr_1][1], cam_mem_add[addr_0][1]} ==  p[4:0]) begin
                  match_flag_carry_3 = 1'b1;
                  pp1 = {2'b10, p[4:0]};
                  break; // exit the loop once a match is found
              end
          end
      end
      
      if( {cam_mem_add[addr_3][0], cam_mem_add[addr_2][0]} == 2'b11) begin
          for (q = 0; q < 32; q = q + 1) begin  
              if ({cam_mem_add[addr_1][0], cam_mem_add[addr_3][1], cam_mem_add[addr_2][1], cam_mem_add[addr_1][1], cam_mem_add[addr_0][1]} ==  q[4:0]) begin
                  match_flag_carry_4 = 1'b1;
                  pp1 = {2'b11, q[4:0]};
                  break; // exit the loop once a match is found
              end
          end
      end
    

  end 
 end
 

  
  assign actual_sum = a+b+c;
  assign sum = {cam_mem[pp1],cam_mem_add[addr_0][0] };
         
endmodule

module adder_64bit_re(
input bit clk,
input  logic rst, 
  input logic write_en,
  input logic [63:0] a, b,c,
  input logic [2:0] data_add [63:0],
  input logic [4:0] data [127:0],
  output logic [64:0] sum, actual_sum,
  output logic [12:0] final_flag
    );
logic [12:0] address0, address1, address2, address3, address4, address5, 
                 address6, address7, address8, address9, address10;
logic [4:0] sub_sum_0, sub_actual_sum_0;
logic [4:0] sub_sum_1, sub_actual_sum_1;
  logic [4:0] sub_sum_2, sub_actual_sum_2;
  logic [4:0] sub_sum_3, sub_actual_sum_3;
  logic [4:0] sub_sum_4, sub_actual_sum_4;
  logic [4:0] sub_sum_5, sub_actual_sum_5;
  logic [4:0] sub_sum_6, sub_actual_sum_6;
  logic [4:0] sub_sum_7, sub_actual_sum_7;
  logic [4:0] sub_sum_8, sub_actual_sum_8;
  logic [4:0] sub_sum_9, sub_actual_sum_9;
  logic [4:0] sub_sum_10, sub_actual_sum_10;
  logic [4:0] sub_sum_11, sub_actual_sum_11;
  logic [4:0] sub_sum_12, sub_actual_sum_12;
  logic [4:0] sub_sum_13, sub_actual_sum_13;
  logic [4:0] sub_sum_14, sub_actual_sum_14;
  logic [4:0] sub_sum_15, sub_actual_sum_15;
  logic [4:0] sub_sum_16, sub_actual_sum_16;
  logic [4:0] sub_sum_17, sub_actual_sum_17;
  logic final_flag0,final_flag1,final_flag2,final_flag3,final_flag4,final_flag5,final_flag6,final_flag7,final_flag8,final_flag9;
  logic final_flag10,final_flag11,final_flag12,final_flag13,final_flag14,final_flag15,final_flag16,final_flag17;
  
logic [32:0] sum_temp,sum_temp0,sum_temp1,sum_temp2,sum_temp3,sum_temp4;
    
  adder_4bit_re add32_0(clk, 1'b1, a[3:0],   b[3:0],   4'b0, data_add, data, sub_sum_0, sub_actual_sum_0, final_flag0);
adder_4bit_re add32_1(clk, 1'b1, a[7:4],   b[7:4],   {3'b0, sub_sum_0[4]}, data_add, data, sub_sum_1, sub_actual_sum_1, final_flag1);
adder_4bit_re add32_2(clk, 1'b1, a[11:8],  b[11:8],  {3'b0, sub_sum_1[4]}, data_add, data, sub_sum_2, sub_actual_sum_2, final_flag2);
adder_4bit_re add32_3(clk, 1'b1, a[15:12], b[15:12], {3'b0, sub_sum_2[4]}, data_add, data, sub_sum_3, sub_actual_sum_3, final_flag3);
adder_4bit_re add32_4(clk, 1'b1, a[19:16], b[19:16], {3'b0, sub_sum_3[4]}, data_add, data, sub_sum_4, sub_actual_sum_4, final_flag4);
adder_4bit_re add32_5(clk, 1'b1, a[23:20], b[23:20], {3'b0, sub_sum_4[4]}, data_add, data, sub_sum_5, sub_actual_sum_5, final_flag5);
adder_4bit_re add32_6(clk, 1'b1, a[27:24], b[27:24], {3'b0, sub_sum_5[4]}, data_add, data, sub_sum_6, sub_actual_sum_6, final_flag6);
adder_4bit_re add32_7(clk, 1'b1, a[31:28], b[31:28], {3'b0, sub_sum_6[4]}, data_add, data, sub_sum_7, sub_actual_sum_7, final_flag7); 
adder_4bit_re add32_8(clk, 1'b1, a[35:32], b[35:32], {3'b0, sub_sum_7[4]}, data_add, data, sub_sum_8, sub_actual_sum_8, final_flag8);
adder_4bit_re add32_9(clk, 1'b1, a[39:36], b[39:36], {3'b0, sub_sum_8[4]}, data_add, data, sub_sum_9, sub_actual_sum_9, final_flag9);
adder_4bit_re add32_10(clk, 1'b1, a[43:40], b[43:40], {3'b0, sub_sum_9[4]}, data_add, data, sub_sum_10, sub_actual_sum_10, final_flag10);
adder_4bit_re add32_11(clk, 1'b1, a[47:44], b[47:44], {3'b0, sub_sum_10[4]}, data_add, data, sub_sum_11, sub_actual_sum_11, final_flag11);
adder_4bit_re add32_12(clk, 1'b1, a[51:48], b[51:48], {3'b0, sub_sum_11[4]}, data_add, data, sub_sum_12, sub_actual_sum_12, final_flag12);
adder_4bit_re add32_13(clk, 1'b1, a[55:52], b[55:52], {3'b0, sub_sum_12[4]}, data_add, data, sub_sum_13, sub_actual_sum_13, final_flag13);
adder_4bit_re add32_14(clk, 1'b1, a[59:56], b[59:56], {3'b0, sub_sum_13[4]}, data_add, data, sub_sum_14, sub_actual_sum_14, final_flag14);
adder_4bit_re add32_15(clk, 1'b1, a[63:60], b[63:60], {3'b0, sub_sum_14[4]}, data_add, data, sub_sum_15, sub_actual_sum_15, final_flag15);

    
assign actual_sum = a+b;
assign final_flag = final_flag7;
always_comb begin
 sum_temp =a+b+c;

end

assign sum = { sub_sum_15, sub_sum_14[3:0], 
              sub_sum_13[3:0], sub_sum_12[3:0], sub_sum_11[3:0], sub_sum_10[3:0], 
              sub_sum_9[3:0], sub_sum_8[3:0], sub_sum_7[3:0], sub_sum_6[3:0], 
              sub_sum_5[3:0], sub_sum_4[3:0], sub_sum_3[3:0], sub_sum_2[3:0], 
              sub_sum_1[3:0], sub_sum_0[3:0]};

/*
  ff sai0(clk,rst,sum_temp,sum_temp0);
   ff sai1(clk,rst,sum_temp0,sum_temp1);
     ff sai2(clk,rst,sum_temp1,sum_temp2);
       ff sai3(clk,rst,sum_temp2,sum_temp3); 
      //   ff sai4(clk,rst,sum_temp3,sum_temp4);

 always_comb begin
actual_sum =sum_temp3;
  
 end

assign sum = {sub_sum_7,sub_sum_6[3:0], sub_sum_5[3:0], sub_sum_4[3:0], sub_sum_3[3:0],sub_sum_2[3:0], sub_sum_1[3:0], sub_sum_0[3:0]};
*/
endmodule


////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module adder_68bit_re(
input bit clk,
input  logic rst, 
  input logic write_en,
  input logic [67:0] a, b,c,
  input logic [2:0] data_add [63:0],
  input logic [4:0] data [127:0],
  output logic [68:0] sum, actual_sum,
  output logic [12:0] final_flag
    );
logic [12:0] address0, address1, address2, address3, address4, address5, 
                 address6, address7, address8, address9, address10;
logic [4:0] sub_sum_0, sub_actual_sum_0;
logic [4:0] sub_sum_1, sub_actual_sum_1;
  logic [4:0] sub_sum_2, sub_actual_sum_2;
  logic [4:0] sub_sum_3, sub_actual_sum_3;
  logic [4:0] sub_sum_4, sub_actual_sum_4;
  logic [4:0] sub_sum_5, sub_actual_sum_5;
  logic [4:0] sub_sum_6, sub_actual_sum_6;
  logic [4:0] sub_sum_7, sub_actual_sum_7;
  logic [4:0] sub_sum_8, sub_actual_sum_8;
  logic [4:0] sub_sum_9, sub_actual_sum_9;
  logic [4:0] sub_sum_10, sub_actual_sum_10;
  logic [4:0] sub_sum_11, sub_actual_sum_11;
  logic [4:0] sub_sum_12, sub_actual_sum_12;
  logic [4:0] sub_sum_13, sub_actual_sum_13;
  logic [4:0] sub_sum_14, sub_actual_sum_14;
  logic [4:0] sub_sum_15, sub_actual_sum_15;
  logic [4:0] sub_sum_16, sub_actual_sum_16;
  logic [4:0] sub_sum_17, sub_actual_sum_17;
  logic final_flag0,final_flag1,final_flag2,final_flag3,final_flag4,final_flag5,final_flag6,final_flag7,final_flag8,final_flag9;
  logic final_flag10,final_flag11,final_flag12,final_flag13,final_flag14,final_flag15,final_flag16,final_flag17;
  
logic [32:0] sum_temp,sum_temp0,sum_temp1,sum_temp2,sum_temp3,sum_temp4;
    
  adder_4bit_re add32_0(clk, 1'b1, a[3:0],   b[3:0],   4'b0, data_add, data, sub_sum_0, sub_actual_sum_0, final_flag0);
adder_4bit_re add32_1(clk, 1'b1, a[7:4],   b[7:4],   {3'b0, sub_sum_0[4]}, data_add, data, sub_sum_1, sub_actual_sum_1, final_flag1);
adder_4bit_re add32_2(clk, 1'b1, a[11:8],  b[11:8],  {3'b0, sub_sum_1[4]}, data_add, data, sub_sum_2, sub_actual_sum_2, final_flag2);
adder_4bit_re add32_3(clk, 1'b1, a[15:12], b[15:12], {3'b0, sub_sum_2[4]}, data_add, data, sub_sum_3, sub_actual_sum_3, final_flag3);
adder_4bit_re add32_4(clk, 1'b1, a[19:16], b[19:16], {3'b0, sub_sum_3[4]}, data_add, data, sub_sum_4, sub_actual_sum_4, final_flag4);
adder_4bit_re add32_5(clk, 1'b1, a[23:20], b[23:20], {3'b0, sub_sum_4[4]}, data_add, data, sub_sum_5, sub_actual_sum_5, final_flag5);
adder_4bit_re add32_6(clk, 1'b1, a[27:24], b[27:24], {3'b0, sub_sum_5[4]}, data_add, data, sub_sum_6, sub_actual_sum_6, final_flag6);
adder_4bit_re add32_7(clk, 1'b1, a[31:28], b[31:28], {3'b0, sub_sum_6[4]}, data_add, data, sub_sum_7, sub_actual_sum_7, final_flag7); 
adder_4bit_re add32_8(clk, 1'b1, a[35:32], b[35:32], {3'b0, sub_sum_7[4]}, data_add, data, sub_sum_8, sub_actual_sum_8, final_flag8);
adder_4bit_re add32_9(clk, 1'b1, a[39:36], b[39:36], {3'b0, sub_sum_8[4]}, data_add, data, sub_sum_9, sub_actual_sum_9, final_flag9);
adder_4bit_re add32_10(clk, 1'b1, a[43:40], b[43:40], {3'b0, sub_sum_9[4]}, data_add, data, sub_sum_10, sub_actual_sum_10, final_flag10);
adder_4bit_re add32_11(clk, 1'b1, a[47:44], b[47:44], {3'b0, sub_sum_10[4]}, data_add, data, sub_sum_11, sub_actual_sum_11, final_flag11);
adder_4bit_re add32_12(clk, 1'b1, a[51:48], b[51:48], {3'b0, sub_sum_11[4]}, data_add, data, sub_sum_12, sub_actual_sum_12, final_flag12);
adder_4bit_re add32_13(clk, 1'b1, a[55:52], b[55:52], {3'b0, sub_sum_12[4]}, data_add, data, sub_sum_13, sub_actual_sum_13, final_flag13);
adder_4bit_re add32_14(clk, 1'b1, a[59:56], b[59:56], {3'b0, sub_sum_13[4]}, data_add, data, sub_sum_14, sub_actual_sum_14, final_flag14);
adder_4bit_re add32_15(clk, 1'b1, a[63:60], b[63:60], {3'b0, sub_sum_14[4]}, data_add, data, sub_sum_15, sub_actual_sum_15, final_flag15);
adder_4bit_re add32_16(clk, 1'b1, a[67:64], b[67:64], {3'b0, sub_sum_15[4]}, data_add, data, sub_sum_16, sub_actual_sum_16, final_flag16);

    
assign actual_sum = a+b;
assign final_flag = final_flag7;
always_comb begin
 sum_temp =a+b+c;

end

assign sum = { sub_sum_16, sub_sum_15[3:0], sub_sum_14[3:0], 
              sub_sum_13[3:0], sub_sum_12[3:0], sub_sum_11[3:0], sub_sum_10[3:0], 
              sub_sum_9[3:0], sub_sum_8[3:0], sub_sum_7[3:0], sub_sum_6[3:0], 
              sub_sum_5[3:0], sub_sum_4[3:0], sub_sum_3[3:0], sub_sum_2[3:0], 
              sub_sum_1[3:0], sub_sum_0[3:0]};


endmodule

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module adder_72bit_re(
input bit clk,
input  logic rst, 
  input logic write_en,
  input logic [71:0] a, b,c,
  input logic [2:0] data_add [63:0],
  input logic [4:0] data [127:0],
  output logic [72:0] sum, actual_sum,
  output logic [12:0] final_flag
    );
logic [12:0] address0, address1, address2, address3, address4, address5, 
                 address6, address7, address8, address9, address10;
logic [4:0] sub_sum_0, sub_actual_sum_0;
logic [4:0] sub_sum_1, sub_actual_sum_1;
  logic [4:0] sub_sum_2, sub_actual_sum_2;
  logic [4:0] sub_sum_3, sub_actual_sum_3;
  logic [4:0] sub_sum_4, sub_actual_sum_4;
  logic [4:0] sub_sum_5, sub_actual_sum_5;
  logic [4:0] sub_sum_6, sub_actual_sum_6;
  logic [4:0] sub_sum_7, sub_actual_sum_7;
  logic [4:0] sub_sum_8, sub_actual_sum_8;
  logic [4:0] sub_sum_9, sub_actual_sum_9;
  logic [4:0] sub_sum_10, sub_actual_sum_10;
  logic [4:0] sub_sum_11, sub_actual_sum_11;
  logic [4:0] sub_sum_12, sub_actual_sum_12;
  logic [4:0] sub_sum_13, sub_actual_sum_13;
  logic [4:0] sub_sum_14, sub_actual_sum_14;
  logic [4:0] sub_sum_15, sub_actual_sum_15;
  logic [4:0] sub_sum_16, sub_actual_sum_16;
  logic [4:0] sub_sum_17, sub_actual_sum_17;
  logic final_flag0,final_flag1,final_flag2,final_flag3,final_flag4,final_flag5,final_flag6,final_flag7,final_flag8,final_flag9;
  logic final_flag10,final_flag11,final_flag12,final_flag13,final_flag14,final_flag15,final_flag16,final_flag17;
  
logic [32:0] sum_temp,sum_temp0,sum_temp1,sum_temp2,sum_temp3,sum_temp4;
    
  adder_4bit_re add32_0(clk, 1'b1, a[3:0],   b[3:0],   4'b0, data_add, data, sub_sum_0, sub_actual_sum_0, final_flag0);
  adder_4bit_re add32_1(clk, 1'b1, a[7:4],   b[7:4],   {3'b0, sub_sum_0[4]}, data_add, data, sub_sum_1, sub_actual_sum_1, final_flag1);
  adder_4bit_re add32_2(clk, 1'b1, a[11:8],  b[11:8],  {3'b0, sub_sum_1[4]}, data_add, data, sub_sum_2, sub_actual_sum_2, final_flag2);
  adder_4bit_re add32_3(clk, 1'b1, a[15:12], b[15:12], {3'b0, sub_sum_2[4]}, data_add, data, sub_sum_3, sub_actual_sum_3, final_flag3);
  adder_4bit_re add32_4(clk, 1'b1, a[19:16], b[19:16], {3'b0, sub_sum_3[4]}, data_add, data, sub_sum_4, sub_actual_sum_4, final_flag4);
  adder_4bit_re add32_5(clk, 1'b1, a[23:20], b[23:20], {3'b0, sub_sum_4[4]}, data_add, data, sub_sum_5, sub_actual_sum_5, final_flag5);
  adder_4bit_re add32_6(clk, 1'b1, a[27:24], b[27:24], {3'b0, sub_sum_5[4]}, data_add, data, sub_sum_6, sub_actual_sum_6, final_flag6);
  adder_4bit_re add32_7(clk, 1'b1, a[31:28], b[31:28], {3'b0, sub_sum_6[4]}, data_add, data, sub_sum_7, sub_actual_sum_7, final_flag7); 
  adder_4bit_re add32_8(clk, 1'b1, a[35:32], b[35:32], {3'b0, sub_sum_7[4]}, data_add, data, sub_sum_8, sub_actual_sum_8, final_flag8);
  adder_4bit_re add32_9(clk, 1'b1, a[39:36], b[39:36], {3'b0, sub_sum_8[4]}, data_add, data, sub_sum_9, sub_actual_sum_9, final_flag9);
  adder_4bit_re add32_10(clk, 1'b1, a[43:40], b[43:40], {3'b0, sub_sum_9[4]}, data_add, data, sub_sum_10, sub_actual_sum_10, final_flag10);
  adder_4bit_re add32_11(clk, 1'b1, a[47:44], b[47:44], {3'b0, sub_sum_10[4]}, data_add, data, sub_sum_11, sub_actual_sum_11, final_flag11);
  adder_4bit_re add32_12(clk, 1'b1, a[51:48], b[51:48], {3'b0, sub_sum_11[4]}, data_add, data, sub_sum_12, sub_actual_sum_12, final_flag12);
  adder_4bit_re add32_13(clk, 1'b1, a[55:52], b[55:52], {3'b0, sub_sum_12[4]}, data_add, data, sub_sum_13, sub_actual_sum_13, final_flag13);
  adder_4bit_re add32_14(clk, 1'b1, a[59:56], b[59:56], {3'b0, sub_sum_13[4]}, data_add, data, sub_sum_14, sub_actual_sum_14, final_flag14);
  adder_4bit_re add32_15(clk, 1'b1, a[63:60], b[63:60], {3'b0, sub_sum_14[4]}, data_add, data, sub_sum_15, sub_actual_sum_15, final_flag15);
  adder_4bit_re add32_16(clk, 1'b1, a[67:64], b[67:64], {3'b0, sub_sum_15[4]}, data_add, data, sub_sum_16, sub_actual_sum_16, final_flag16);
  adder_4bit_re add32_17(clk, 1'b1, a[71:68], b[71:68], {3'b0, sub_sum_16[4]}, data_add, data, sub_sum_17, sub_actual_sum_17, final_flag17);


    
assign actual_sum = a+b;
assign final_flag = final_flag7;
always_comb begin
 sum_temp =a+b+c;

end

assign sum = { sub_sum_17,sub_sum_16[3:0], sub_sum_15[3:0], sub_sum_14[3:0], 
              sub_sum_13[3:0], sub_sum_12[3:0], sub_sum_11[3:0], sub_sum_10[3:0], 
              sub_sum_9[3:0], sub_sum_8[3:0], sub_sum_7[3:0], sub_sum_6[3:0], 
              sub_sum_5[3:0], sub_sum_4[3:0], sub_sum_3[3:0], sub_sum_2[3:0], 
              sub_sum_1[3:0], sub_sum_0[3:0]};


endmodule











///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// count ones in coloum of 7 length
//seems no chnages requried || change in data
module count_ones_sub(
input logic a,b,c,d,e,f,
input logic [2:0] data [63:0],
output logic [2:0] sub_out // 3 bit output 1+1+1+1+1+1= 110
    );

  logic [2:0] sub_out0,sub_out1,sub_out2; // 3 bit output 1+1+1+1 = 100
  logic out0_flag,out1_flag,out2_flag;
  logic [2:0] add [63:0];
  int j,k,l,u;
  logic [3:0] sub_sum;
  logic data_flag;
  logic [3:0] sub_out_actual;
  assign sub_out_actual = a+b+c+d+e+f;
  
  
    always_comb begin 
    for (u = 0; u< 64; u++) begin
      add[u] = data[u];  // Only assign the lower 2 bits to `add`
    end
    data_flag = 1'b1;
  end

always_comb begin 
sub_out0 = 2'b0;
out0_flag = 1'b0;
if (data_flag) begin
  for(l=0; l<64;l++) begin
    if({a,b,c,d,e,f} == l[5:0]) begin
      sub_out0 = add[l[5:0]]; // add[111111]
      out0_flag = 1'b1;
  break;
end
end
end
end

assign sub_out = sub_out0;

endmodule


///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//8 cycles
module count_mul_v2(
input logic p0, p1, p2, p3, p4, p5, p6, p7, p8, p9, p10, p11, p12, p13, p14, p15, p16, p17, p18, p19, p20, p21, p22, p23, p24, p25, p26, p27, p28, p29, p30, p31,
input logic [2:0] data [63:0],
input logic [4:0] data_unq [127:0],
input logic clk,
output logic [5:0] out //7 bit output becaus 32 x1  = 32 
    );
    
  logic [2:0] out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10,out11,out12; // adding 5 single bits  = 3 bit output
  logic out0_flag, out1_flag, out2_flag, out3_flag, out4_flag, out5_flag, out6_flag, out7_flag, out8_flag, out9_flag, out10_flag,out11_flag,out12_flag;
  logic [2:0] add [63:0];
  int loop_0, loop_1, loop_2, loop_3, loop_4, loop_5, loop_6, loop_7, loop_8, loop_9, loop_10,loop_11,loop_12,loop_data,loop_data1;
  logic [5:0] sum;
  logic [5:0] actual_sum_v2;
  logic [2:0] sum0,sum1,sum2;
  logic data_flag,data_flag1;

   logic [12:0] address_v2;
   logic  [4:0] cam_mem_unq [127:0]; // CAM cell 
  
  
  
   always_ff @(posedge clk) begin 
    for (loop_data = 0; loop_data< 64; loop_data++) begin
      add[loop_data] = data[loop_data];  // Only assign the lower 2 bits to `add`
    end
    data_flag1 = 1'b1;
  end
    
   always_ff @(posedge clk) begin 
    for (loop_data1 = 0; loop_data1< 128; loop_data1++) begin
      cam_mem_unq[loop_data1] = data_unq[loop_data1];  // Only assign the lower 2 bits to `add`
    end
    data_flag = 1'b1;
  end

  

 always_ff @(posedge clk) begin
  out0 = 3'b0;
    out0_flag = 1'b0;
    if (data_flag) begin
     for(loop_0=0; loop_0<64;loop_0++) begin
        if({p0,p1,p2,p3,p4,p5} == loop_0[5:0]) begin
     out0 = add[loop_0[5:0]];
      out0_flag = 1'b1;
      break;
    end
  end
  end
end
 always_ff @(posedge clk) begin
  out1 = 3'b0;
    out1_flag = 1'b0;
    if (data_flag) begin
     for(loop_1=0; loop_1<64;loop_1++) begin
        if({p6,p7,p8,p9,p10,p11} == loop_1[5:0]) begin
     out1 = add[loop_1[5:0]];
      out1_flag = 1'b1;
      break;
    end
  end
  end
end
 always_ff @(posedge clk) begin
  out2 = 3'b0;
    out2_flag = 1'b0;
    if (data_flag) begin
     for(loop_2=0; loop_2<64;loop_2++) begin
        if({p12,p13,p14,p15,p16,p17} == loop_2[5:0]) begin
     out2 = add[loop_2[5:0]];
      out2_flag = 1'b1;
      break;
    end
  end
  end
end
 always_ff @(posedge clk) begin
  out3 = 3'b0;
    out3_flag = 1'b0;
    if (data_flag) begin
     for(loop_3=0; loop_3<64;loop_3++) begin
        if({p18,p19,p20,p21,p22,p23} == loop_3[5:0]) begin
     out3 = add[loop_3[5:0]];
      out3_flag = 1'b1;
      break;
    end
  end
  end
end
 always_ff @(posedge clk) begin
  out4 = 3'b0;
    out4_flag = 1'b0;
    if (data_flag) begin
     for(loop_4=0; loop_4<64;loop_4++) begin
        if({p24,p25,p26,p27,p28,p29} == loop_4[5:0]) begin
     out4 = add[loop_4[5:0]];
      out4_flag = 1'b1;
      break;
    end
  end
  end
end
 always_ff @(posedge clk) begin
  out5 = 3'b0;
    out5_flag = 1'b0;
    if (data_flag) begin
     for(loop_5=0; loop_5<64;loop_5++) begin
        if({1'b0,1'b0,1'b0,1'b0,p30,p31} == loop_5[5:0]) begin
     out5 = add[loop_5[5:0]];
      out5_flag = 1'b1;
      break;
    end
  end
  end
end

//////////////////////////////////////////////////////////////////////////////////////////
// count the all 7 3bit number columns
//////////////////////////////////////////////////////////////////////////////////////////
count_ones_sub sub0(
    .a(out0[0]),
    .b(out1[0]),
    .c(out2[0]),
    .d(out3[0]),
    .e(out4[0]),
    .f(out5[0]),
    .data(add),
    .sub_out(sum0)
);

count_ones_sub sub1(
    .a(out0[1]),
    .b(out1[1]),
    .c(out2[1]),
    .d(out3[1]),
    .e(out4[1]),
    .f(out5[1]),
    .data(add),
    .sub_out(sum1)
);

count_ones_sub sub2(
    .a(out0[2]),
    .b(out1[2]),
    .c(out2[2]),
    .d(out3[2]),
    .e(out4[2]),
    .f(out5[2]),
    .data(add),
    .sub_out(sum2)
);

 

  adder_4bit_re s1(
    .clk(clk),
    .write_en(1'b1),
    .a({1'b0,1'b0,sum0[2:1]}),
    .b({1'b0,sum1}),
    .c({sum2,1'b0}),
    .data_add(add),
    .data_unq(cam_mem_unq),
    .sum(sum),
    .actual_sum(actual_sum_v2),
    .address(address_v2)
  );

assign out = {sum,sum0[0]};

endmodule


module adder_mul_64bit_re(
input logic clk,
input logic rst,
  input logic write_en,
  input logic [63:0] p0, p1, p2, p3, p4, p5, p6, p7, p8, p9, p10, p11, p12, p13, p14, p15,
        p16, p17, p18, p19, p20, p21, p22, p23, p24, p25, p26, p27, p28, p29, p30, p31,
  input logic  [2:0] data [63:0],
  input logic [4:0] data_unq [127:0],
  output logic [72:0] sum, actual_sum,
  output logic [12:0] address

    );
   
   logic [72:0] actualsum_pps, actualsum_pps01_23_45;
   logic [64:0] sum_pps45,sum_pps23,sum_pps01;
    logic [64:0] actual_sum23,actual_sum01,actual_sum45;
    
      logic [68:0]  actual_sum0123,sum_pps0123;
      logic [72:0] sum_pps012345,actual_sum012345;

   
   logic [5:0] count0, count1, count2, count3, count4, count5, count6, count7, 
                count8, count9, count10, count11, count12, count13, count14, count15,
                count16, count17, count18, count19, count20, count21, 
                count22, count23, count24, count25, count26,count27, count28, count29, count30, 
                count31, count32, count33, count34, count35, count36, count37, count38, count39, 
                count40, count41, count42, count43, count44, count45, count46, count47, count48, 
                count49, count50, count51, count52, count53, count54, count55, count56, count57, 
                count58, count59, count60, count61, count62, count63;
   
                


logic final_flag,final_flag01,final_flag23,final_flag45,final_flag012345,final_flag0123;
logic [68:0] pps0, pps1, pps2, pps3,pps4,pps5;



    
 assign actual_sum =p0 + p1 + p2 + p3 + p4 + p5 + p6 + p7 + p8 + p9 + p10 + p11 + p12 + p13 + p14 + p15 + p16 + p17 + p18 + p19 + p20 + p21 + p22 + p23 + p24 + p25 + p26 + p27 + p28 + p29 + p30 + p31;
   
count_mul_v2 x10(p0[0], p1[0], p2[0], p3[0], p4[0], p5[0], p6[0], p7[0], p8[0], p9[0], p10[0], p11[0], p12[0], p13[0], p14[0], p15[0], p16[0], p17[0], p18[0], p19[0], p20[0], p21[0], p22[0], p23[0], p24[0], p25[0], p26[0], p27[0],  p28[0], p29[0], p30[0], p31[0], data,data_unq,clk, count0); 
 count_mul_v2 x11(p0[1], p1[1], p2[1], p3[1], p4[1], p5[1], p6[1], p7[1], p8[1], p9[1], p10[1], p11[1], p12[1], p13[1], p14[1], p15[1], p16[1], p17[1], p18[1], p19[1], p20[1], p21[1], p22[1], p23[1], p24[1], p25[1], p26[1], p27[1], 
 p28[1], p29[1], p30[1], p31[1], data,data_unq,clk, count1); 
 count_mul_v2 x12(p0[2], p1[2], p2[2], p3[2], p4[2], p5[2], p6[2], p7[2], p8[2], p9[2], p10[2], p11[2], p12[2], p13[2], p14[2], p15[2], p16[2], p17[2], p18[2], p19[2], p20[2], p21[2], p22[2], p23[2], p24[2], p25[2], p26[2], p27[2], 
 p28[2], p29[2], p30[2], p31[2], data,data_unq,clk, count2); 
 count_mul_v2 x13(p0[3], p1[3], p2[3], p3[3], p4[3], p5[3], p6[3], p7[3], p8[3], p9[3], p10[3], p11[3], p12[3], p13[3], p14[3], p15[3], p16[3], p17[3], p18[3], p19[3], p20[3], p21[3], p22[3], p23[3], p24[3], p25[3], p26[3], p27[3], 
 p28[3], p29[3], p30[3], p31[3], data,data_unq,clk, count3); 
 count_mul_v2 x14(p0[4], p1[4], p2[4], p3[4], p4[4], p5[4], p6[4], p7[4], p8[4], p9[4], p10[4], p11[4], p12[4], p13[4], p14[4], p15[4], p16[4], p17[4], p18[4], p19[4], p20[4], p21[4], p22[4], p23[4], p24[4], p25[4], p26[4], p27[4], 
 p28[4], p29[4], p30[4], p31[4], data,data_unq,clk, count4); 
 count_mul_v2 x15(p0[5], p1[5], p2[5], p3[5], p4[5], p5[5], p6[5], p7[5], p8[5], p9[5], p10[5], p11[5], p12[5], p13[5], p14[5], p15[5], p16[5], p17[5], p18[5], p19[5], p20[5], p21[5], p22[5], p23[5], p24[5], p25[5], p26[5], p27[5], 
 p28[5], p29[5], p30[5], p31[5], data,data_unq,clk, count5); 
 count_mul_v2 x16(p0[6], p1[6], p2[6], p3[6], p4[6], p5[6], p6[6], p7[6], p8[6], p9[6], p10[6], p11[6], p12[6], p13[6], p14[6], p15[6], p16[6], p17[6], p18[6], p19[6], p20[6], p21[6], p22[6], p23[6], p24[6], p25[6], p26[6], p27[6], 
 p28[6], p29[6], p30[6], p31[6], data,data_unq,clk, count6); 
 count_mul_v2 x17(p0[7], p1[7], p2[7], p3[7], p4[7], p5[7], p6[7], p7[7], p8[7], p9[7], p10[7], p11[7], p12[7], p13[7], p14[7], p15[7], p16[7], p17[7], p18[7], p19[7], p20[7], p21[7], p22[7], p23[7], p24[7], p25[7], p26[7], p27[7], 
 p28[7], p29[7], p30[7], p31[7], data,data_unq,clk, count7); 
 count_mul_v2 x18(p0[8], p1[8], p2[8], p3[8], p4[8], p5[8], p6[8], p7[8], p8[8], p9[8], p10[8], p11[8], p12[8], p13[8], p14[8], p15[8], p16[8], p17[8], p18[8], p19[8], p20[8], p21[8], p22[8], p23[8], p24[8], p25[8], p26[8], p27[8], 
 p28[8], p29[8], p30[8], p31[8], data,data_unq,clk, count8); 
 count_mul_v2 x19(p0[9], p1[9], p2[9], p3[9], p4[9], p5[9], p6[9], p7[9], p8[9], p9[9], p10[9], p11[9], p12[9], p13[9], p14[9], p15[9], p16[9], p17[9], p18[9], p19[9], p20[9], p21[9], p22[9], p23[9], p24[9], p25[9], p26[9], p27[9], 
 p28[9], p29[9], p30[9], p31[9], data,data_unq,clk, count9); 
 count_mul_v2 x20(p0[10], p1[10], p2[10], p3[10], p4[10], p5[10], p6[10], p7[10], p8[10], p9[10], p10[10], p11[10], p12[10], p13[10], p14[10], p15[10], p16[10], p17[10], p18[10], p19[10], p20[10], p21[10], p22[10], p23[10], p24[10], p25[10], p26[10], p27[10], p28[10], p29[10], p30[10], p31[10], data,data_unq,clk, count10); 
 count_mul_v2 x21(p0[11], p1[11], p2[11], p3[11], p4[11], p5[11], p6[11], p7[11], p8[11], p9[11], p10[11], p11[11], p12[11], p13[11], p14[11], p15[11], p16[11], p17[11], p18[11], p19[11], p20[11], p21[11], p22[11], p23[11], p24[11], p25[11], p26[11], p27[11], p28[11], p29[11], p30[11], p31[11], data,data_unq,clk, count11); 
 count_mul_v2 x22(p0[12], p1[12], p2[12], p3[12], p4[12], p5[12], p6[12], p7[12], p8[12], p9[12], p10[12], p11[12], p12[12], p13[12], p14[12], p15[12], p16[12], p17[12], p18[12], p19[12], p20[12], p21[12], p22[12], p23[12], p24[12], p25[12], p26[12], p27[12], p28[12], p29[12], p30[12], p31[12], data,data_unq,clk, count12);
 count_mul_v2 x23(p0[13], p1[13], p2[13], p3[13], p4[13], p5[13], p6[13], p7[13], p8[13], p9[13], p10[13], p11[13], p12[13], p13[13], p14[13], p15[13], p16[13], p17[13], p18[13], p19[13], p20[13], p21[13], p22[13], p23[13], p24[13], p25[13], p26[13], p27[13], p28[13], p29[13], p30[13], p31[13], data,data_unq,clk, count13);
 count_mul_v2 x24(p0[14], p1[14], p2[14], p3[14], p4[14], p5[14], p6[14], p7[14], p8[14], p9[14], p10[14], p11[14], p12[14], p13[14], p14[14], p15[14], p16[14], p17[14], p18[14], p19[14], p20[14], p21[14], p22[14], p23[14], p24[14], p25[14], p26[14], p27[14], p28[14], p29[14], p30[14], p31[14], data,data_unq,clk, count14);
 count_mul_v2 x25(p0[15], p1[15], p2[15], p3[15], p4[15], p5[15], p6[15], p7[15], p8[15], p9[15], p10[15], p11[15], p12[15], p13[15], p14[15], p15[15], p16[15], p17[15], p18[15], p19[15], p20[15], p21[15], p22[15], p23[15], p24[15], p25[15], p26[15], p27[15], p28[15], p29[15], p30[15], p31[15], data,data_unq,clk, count15);
 count_mul_v2 x26(p0[16], p1[16], p2[16], p3[16], p4[16], p5[16], p6[16], p7[16], p8[16], p9[16], p10[16], p11[16], p12[16], p13[16], p14[16], p15[16], p16[16], p17[16], p18[16], p19[16], p20[16], p21[16], p22[16], p23[16], p24[16], p25[16], p26[16], p27[16], p28[16], p29[16], p30[16], p31[16], data,data_unq,clk, count16);
 count_mul_v2 x27(p0[17], p1[17], p2[17], p3[17], p4[17], p5[17], p6[17], p7[17], p8[17], p9[17], p10[17], p11[17], p12[17], p13[17], p14[17], p15[17], p16[17], p17[17], p18[17], p19[17], p20[17], p21[17], p22[17], p23[17], p24[17], p25[17], p26[17], p27[17], p28[17], p29[17], p30[17], p31[17], data,data_unq,clk, count17);
 count_mul_v2 x28(p0[18], p1[18], p2[18], p3[18], p4[18], p5[18], p6[18], p7[18], p8[18], p9[18], p10[18], p11[18], p12[18], p13[18], p14[18], p15[18], p16[18], p17[18], p18[18], p19[18], p20[18], p21[18], p22[18], p23[18], p24[18], p25[18], p26[18], p27[18], p28[18], p29[18], p30[18], p31[18], data,data_unq,clk, count18);
 count_mul_v2 x29(p0[19], p1[19], p2[19], p3[19], p4[19], p5[19], p6[19], p7[19], p8[19], p9[19], p10[19], p11[19], p12[19], p13[19], p14[19], p15[19], p16[19], p17[19], p18[19], p19[19], p20[19], p21[19], p22[19], p23[19], p24[19], p25[19], p26[19], p27[19], p28[19], p29[19], p30[19], p31[19], data,data_unq,clk, count19);
 count_mul_v2 x30(p0[20], p1[20], p2[20], p3[20], p4[20], p5[20], p6[20], p7[20], p8[20], p9[20], p10[20], p11[20], p12[20], p13[20], p14[20], p15[20], p16[20], p17[20], p18[20], p19[20], p20[20], p21[20], p22[20], p23[20], p24[20], p25[20], p26[20], p27[20], p28[20], p29[20], p30[20], p31[20], data,data_unq,clk, count20);
 count_mul_v2 x31(p0[21], p1[21], p2[21], p3[21], p4[21], p5[21], p6[21], p7[21], p8[21], p9[21], p10[21], p11[21], p12[21], p13[21], p14[21], p15[21], p16[21], p17[21], p18[21], p19[21], p20[21], p21[21], p22[21], p23[21], p24[21], p25[21], p26[21], p27[21], p28[21], p29[21], p30[21], p31[21], data,data_unq,clk, count21);
 count_mul_v2 x32(p0[22], p1[22], p2[22], p3[22], p4[22], p5[22], p6[22], p7[22], p8[22], p9[22], p10[22], p11[22], p12[22], p13[22], p14[22], p15[22], p16[22], p17[22], p18[22], p19[22], p20[22], p21[22], p22[22], p23[22], p24[22], p25[22], p26[22], p27[22], p28[22], p29[22], p30[22], p31[22], data,data_unq,clk, count22);
 count_mul_v2 x33(p0[23], p1[23], p2[23], p3[23], p4[23], p5[23], p6[23], p7[23], p8[23], p9[23], p10[23], p11[23], p12[23], p13[23], p14[23], p15[23], p16[23], p17[23], p18[23], p19[23], p20[23], p21[23], p22[23], p23[23], p24[23], p25[23], p26[23], p27[23], p28[23], p29[23], p30[23], p31[23], data,data_unq,clk, count23);
 count_mul_v2 x34(p0[24], p1[24], p2[24], p3[24], p4[24], p5[24], p6[24], p7[24], p8[24], p9[24], p10[24], p11[24], p12[24], p13[24], p14[24], p15[24], p16[24], p17[24], p18[24], p19[24], p20[24], p21[24], p22[24], p23[24], p24[24], p25[24], p26[24], p27[24], p28[24], p29[24], p30[24], p31[24], data,data_unq,clk, count24);
 count_mul_v2 x35(p0[25], p1[25], p2[25], p3[25], p4[25], p5[25], p6[25], p7[25], p8[25], p9[25], p10[25], p11[25], p12[25], p13[25], p14[25], p15[25], p16[25], p17[25], p18[25], p19[25], p20[25], p21[25], p22[25], p23[25], p24[25], p25[25], p26[25], p27[25], p28[25], p29[25], p30[25], p31[25], data,data_unq,clk, count25);
 count_mul_v2 x36(p0[26], p1[26], p2[26], p3[26], p4[26], p5[26], p6[26], p7[26], p8[26], p9[26], p10[26], p11[26], p12[26], p13[26], p14[26], p15[26], p16[26], p17[26], p18[26], p19[26], p20[26], p21[26], p22[26], p23[26], p24[26], p25[26], p26[26], p27[26], p28[26], p29[26], p30[26], p31[26], data,data_unq,clk, count26);
 count_mul_v2 x37(p0[27], p1[27], p2[27], p3[27], p4[27], p5[27], p6[27], p7[27], p8[27], p9[27], p10[27], p11[27], p12[27], p13[27], p14[27], p15[27], p16[27], p17[27], p18[27], p19[27], p20[27], p21[27], p22[27], p23[27], p24[27], p25[27], p26[27], p27[27], p28[27], p29[27], p30[27], p31[27], data,data_unq,clk, count27);
 count_mul_v2 x38(p0[28], p1[28], p2[28], p3[28], p4[28], p5[28], p6[28], p7[28], p8[28], p9[28], p10[28], p11[28], p12[28], p13[28], p14[28], p15[28], p16[28], p17[28], p18[28], p19[28], p20[28], p21[28], p22[28], p23[28], p24[28], p25[28], p26[28], p27[28], p28[28], p29[28], p30[28], p31[28], data,data_unq,clk, count28);
 count_mul_v2 x39(p0[29], p1[29], p2[29], p3[29], p4[29], p5[29], p6[29], p7[29], p8[29], p9[29], p10[29], p11[29], p12[29], p13[29], p14[29], p15[29], p16[29], p17[29], p18[29], p19[29], p20[29], p21[29], p22[29], p23[29], p24[29], p25[29], p26[29], p27[29], p28[29], p29[29], p30[29], p31[29], data,data_unq,clk, count29);
 count_mul_v2 x40(p0[30], p1[30], p2[30], p3[30], p4[30], p5[30], p6[30], p7[30], p8[30], p9[30], p10[30], p11[30], p12[30], p13[30], p14[30], p15[30], p16[30], p17[30], p18[30], p19[30], p20[30], p21[30], p22[30], p23[30], p24[30], p25[30], p26[30], p27[30], p28[30], p29[30], p30[30], p31[30], data,data_unq,clk, count30);
 count_mul_v2 x41(p0[31], p1[31], p2[31], p3[31], p4[31], p5[31], p6[31], p7[31], p8[31], p9[31], p10[31], p11[31], p12[31], p13[31], p14[31], p15[31], p16[31], p17[31], p18[31], p19[31], p20[31], p21[31], p22[31], p23[31], p24[31], p25[31], p26[31], p27[31], p28[31], p29[31], p30[31], p31[31], data,data_unq,clk, count31);
 count_mul_v2 x42(p0[32], p1[32], p2[32], p3[32], p4[32], p5[32], p6[32], p7[32], p8[32], p9[32], p10[32], p11[32], p12[32], p13[32], p14[32], p15[32], p16[32], p17[32], p18[32], p19[32], p20[32], p21[32], p22[32], p23[32], p24[32], p25[32], p26[32], p27[32], p28[32], p29[32], p30[32], p31[32], data,data_unq,clk, count32);
 count_mul_v2 x43(p0[33], p1[33], p2[33], p3[33], p4[33], p5[33], p6[33], p7[33], p8[33], p9[33], p10[33], p11[33], p12[33], p13[33], p14[33], p15[33], p16[33], p17[33], p18[33], p19[33], p20[33], p21[33], p22[33], p23[33], p24[33], p25[33], p26[33], p27[33], p28[33], p29[33], p30[33], p31[33], data,data_unq,clk, count33);
 count_mul_v2 x44(p0[34], p1[34], p2[34], p3[34], p4[34], p5[34], p6[34], p7[34], p8[34], p9[34], p10[34], p11[34], p12[34], p13[34], p14[34], p15[34], p16[34], p17[34], p18[34], p19[34], p20[34], p21[34], p22[34], p23[34], p24[34], p25[34], p26[34], p27[34], p28[34], p29[34], p30[34], p31[34], data,data_unq,clk, count34);
 count_mul_v2 x45(p0[35], p1[35], p2[35], p3[35], p4[35], p5[35], p6[35], p7[35], p8[35], p9[35], p10[35], p11[35], p12[35], p13[35], p14[35], p15[35], p16[35], p17[35], p18[35], p19[35], p20[35], p21[35], p22[35], p23[35], p24[35], p25[35], p26[35], p27[35], p28[35], p29[35], p30[35], p31[35], data,data_unq,clk, count35);
 count_mul_v2 x46(p0[36], p1[36], p2[36], p3[36], p4[36], p5[36], p6[36], p7[36], p8[36], p9[36], p10[36], p11[36], p12[36], p13[36], p14[36], p15[36], p16[36], p17[36], p18[36], p19[36], p20[36], p21[36], p22[36], p23[36], p24[36], p25[36], p26[36], p27[36], p28[36], p29[36], p30[36], p31[36], data,data_unq,clk, count36);
 count_mul_v2 x47(p0[37], p1[37], p2[37], p3[37], p4[37], p5[37], p6[37], p7[37], p8[37], p9[37], p10[37], p11[37], p12[37], p13[37], p14[37], p15[37], p16[37], p17[37], p18[37], p19[37], p20[37], p21[37], p22[37], p23[37], p24[37], p25[37], p26[37], p27[37], p28[37], p29[37], p30[37], p31[37], data,data_unq,clk, count37);
 count_mul_v2 x48(p0[38], p1[38], p2[38], p3[38], p4[38], p5[38], p6[38], p7[38], p8[38], p9[38], p10[38], p11[38], p12[38], p13[38], p14[38], p15[38], p16[38], p17[38], p18[38], p19[38], p20[38], p21[38], p22[38], p23[38], p24[38], p25[38], p26[38], p27[38], p28[38], p29[38], p30[38], p31[38], data,data_unq,clk, count38);
 count_mul_v2 x49(p0[39], p1[39], p2[39], p3[39], p4[39], p5[39], p6[39], p7[39], p8[39], p9[39], p10[39], p11[39], p12[39], p13[39], p14[39], p15[39], p16[39], p17[39], p18[39], p19[39], p20[39], p21[39], p22[39], p23[39], p24[39], p25[39], p26[39], p27[39], p28[39], p29[39], p30[39], p31[39], data,data_unq,clk, count39);
 count_mul_v2 x50(p0[40], p1[40], p2[40], p3[40], p4[40], p5[40], p6[40], p7[40], p8[40], p9[40], p10[40], p11[40], p12[40], p13[40], p14[40], p15[40], p16[40], p17[40], p18[40], p19[40], p20[40], p21[40], p22[40], p23[40], p24[40], p25[40], p26[40], p27[40], p28[40], p29[40], p30[40], p31[40], data,data_unq,clk, count40);
 count_mul_v2 x51(p0[41], p1[41], p2[41], p3[41], p4[41], p5[41], p6[41], p7[41], p8[41], p9[41], p10[41], p11[41], p12[41], p13[41], p14[41], p15[41], p16[41], p17[41], p18[41], p19[41], p20[41], p21[41], p22[41], p23[41], p24[41], p25[41], p26[41], p27[41], p28[41], p29[41], p30[41], p31[41], data,data_unq,clk, count41);
 count_mul_v2 x52(p0[42], p1[42], p2[42], p3[42], p4[42], p5[42], p6[42], p7[42], p8[42], p9[42], p10[42], p11[42], p12[42], p13[42], p14[42], p15[42], p16[42], p17[42], p18[42], p19[42], p20[42], p21[42], p22[42], p23[42], p24[42], p25[42], p26[42], p27[42], p28[42], p29[42], p30[42], p31[42], data,data_unq,clk, count42);
 count_mul_v2 x53(p0[43], p1[43], p2[43], p3[43], p4[43], p5[43], p6[43], p7[43], p8[43], p9[43], p10[43], p11[43], p12[43], p13[43], p14[43], p15[43], p16[43], p17[43], p18[43], p19[43], p20[43], p21[43], p22[43], p23[43], p24[43], p25[43], p26[43], p27[43], p28[43], p29[43], p30[43], p31[43], data,data_unq,clk, count43);
 count_mul_v2 x54(p0[44], p1[44], p2[44], p3[44], p4[44], p5[44], p6[44], p7[44], p8[44], p9[44], p10[44], p11[44], p12[44], p13[44], p14[44], p15[44], p16[44], p17[44], p18[44], p19[44], p20[44], p21[44], p22[44], p23[44], p24[44], p25[44], p26[44], p27[44], p28[44], p29[44], p30[44], p31[44], data,data_unq,clk, count44);
 count_mul_v2 x55(p0[45], p1[45], p2[45], p3[45], p4[45], p5[45], p6[45], p7[45], p8[45], p9[45], p10[45], p11[45], p12[45], p13[45], p14[45], p15[45], p16[45], p17[45], p18[45], p19[45], p20[45], p21[45], p22[45], p23[45], p24[45], p25[45], p26[45], p27[45], p28[45], p29[45], p30[45], p31[45], data,data_unq,clk, count45);
 count_mul_v2 x56(p0[46], p1[46], p2[46], p3[46], p4[46], p5[46], p6[46], p7[46], p8[46], p9[46], p10[46], p11[46], p12[46], p13[46], p14[46], p15[46], p16[46], p17[46], p18[46], p19[46], p20[46], p21[46], p22[46], p23[46], p24[46], p25[46], p26[46], p27[46], p28[46], p29[46], p30[46], p31[46], data,data_unq,clk, count46);
 count_mul_v2 x57(p0[47], p1[47], p2[47], p3[47], p4[47], p5[47], p6[47], p7[47], p8[47], p9[47], p10[47], p11[47], p12[47], p13[47], p14[47], p15[47], p16[47], p17[47], p18[47], p19[47], p20[47], p21[47], p22[47], p23[47], p24[47], p25[47], p26[47], p27[47], p28[47], p29[47], p30[47], p31[47], data,data_unq,clk, count47);
 count_mul_v2 x58(p0[48], p1[48], p2[48], p3[48], p4[48], p5[48], p6[48], p7[48], p8[48], p9[48], p10[48], p11[48], p12[48], p13[48], p14[48], p15[48], p16[48], p17[48], p18[48], p19[48], p20[48], p21[48], p22[48], p23[48], p24[48], p25[48], p26[48], p27[48], p28[48], p29[48], p30[48], p31[48], data,data_unq,clk, count48);
 count_mul_v2 x59(p0[49], p1[49], p2[49], p3[49], p4[49], p5[49], p6[49], p7[49], p8[49], p9[49], p10[49], p11[49], p12[49], p13[49], p14[49], p15[49], p16[49], p17[49], p18[49], p19[49], p20[49], p21[49], p22[49], p23[49], p24[49], p25[49], p26[49], p27[49], p28[49], p29[49], p30[49], p31[49], data,data_unq,clk, count49);
 count_mul_v2 x60(p0[50], p1[50], p2[50], p3[50], p4[50], p5[50], p6[50], p7[50], p8[50], p9[50], p10[50], p11[50], p12[50], p13[50], p14[50], p15[50], p16[50], p17[50], p18[50], p19[50], p20[50], p21[50], p22[50], p23[50], p24[50], p25[50], p26[50], p27[50], p28[50], p29[50], p30[50], p31[50], data,data_unq,clk, count50);
 count_mul_v2 x61(p0[51], p1[51], p2[51], p3[51], p4[51], p5[51], p6[51], p7[51], p8[51], p9[51], p10[51], p11[51], p12[51], p13[51], p14[51], p15[51], p16[51], p17[51], p18[51], p19[51], p20[51], p21[51], p22[51], p23[51], p24[51], p25[51], p26[51], p27[51], p28[51], p29[51], p30[51], p31[51], data,data_unq,clk, count51);
 count_mul_v2 x62(p0[52], p1[52], p2[52], p3[52], p4[52], p5[52], p6[52], p7[52], p8[52], p9[52], p10[52], p11[52], p12[52], p13[52], p14[52], p15[52], p16[52], p17[52], p18[52], p19[52], p20[52], p21[52], p22[52], p23[52], p24[52], p25[52], p26[52], p27[52], p28[52], p29[52], p30[52], p31[52], data,data_unq,clk, count52);
 count_mul_v2 x63(p0[53], p1[53], p2[53], p3[53], p4[53], p5[53], p6[53], p7[53], p8[53], p9[53], p10[53], p11[53], p12[53], p13[53], p14[53], p15[53], p16[53], p17[53], p18[53], p19[53], p20[53], p21[53], p22[53], p23[53], p24[53], p25[53], p26[53], p27[53], p28[53], p29[53], p30[53], p31[53], data,data_unq,clk, count53);
 count_mul_v2 x64(p0[54], p1[54], p2[54], p3[54], p4[54], p5[54], p6[54], p7[54], p8[54], p9[54], p10[54], p11[54], p12[54], p13[54], p14[54], p15[54], p16[54], p17[54], p18[54], p19[54], p20[54], p21[54], p22[54], p23[54], p24[54], p25[54], p26[54], p27[54], p28[54], p29[54], p30[54], p31[54], data,data_unq,clk, count54);
 count_mul_v2 x65(p0[55], p1[55], p2[55], p3[55], p4[55], p5[55], p6[55], p7[55], p8[55], p9[55], p10[55], p11[55], p12[55], p13[55], p14[55], p15[55], p16[55], p17[55], p18[55], p19[55], p20[55], p21[55], p22[55], p23[55], p24[55], p25[55], p26[55], p27[55], p28[55], p29[55], p30[55], p31[55], data,data_unq,clk, count55);
 count_mul_v2 x66(p0[56], p1[56], p2[56], p3[56], p4[56], p5[56], p6[56], p7[56], p8[56], p9[56], p10[56], p11[56], p12[56], p13[56], p14[56], p15[56], p16[56], p17[56], p18[56], p19[56], p20[56], p21[56], p22[56], p23[56], p24[56], p25[56], p26[56], p27[56], p28[56], p29[56], p30[56], p31[56], data,data_unq,clk, count56);
 count_mul_v2 x67(p0[57], p1[57], p2[57], p3[57], p4[57], p5[57], p6[57], p7[57], p8[57], p9[57], p10[57], p11[57], p12[57], p13[57], p14[57], p15[57], p16[57], p17[57], p18[57], p19[57], p20[57], p21[57], p22[57], p23[57], p24[57], p25[57], p26[57], p27[57], p28[57], p29[57], p30[57], p31[57], data,data_unq,clk, count57);
 count_mul_v2 x68(p0[58], p1[58], p2[58], p3[58], p4[58], p5[58], p6[58], p7[58], p8[58], p9[58], p10[58], p11[58], p12[58], p13[58], p14[58], p15[58], p16[58], p17[58], p18[58], p19[58], p20[58], p21[58], p22[58], p23[58], p24[58], p25[58], p26[58], p27[58], p28[58], p29[58], p30[58], p31[58], data,data_unq,clk, count58);
 count_mul_v2 x69(p0[59], p1[59], p2[59], p3[59], p4[59], p5[59], p6[59], p7[59], p8[59], p9[59], p10[59], p11[59], p12[59], p13[59], p14[59], p15[59], p16[59], p17[59], p18[59], p19[59], p20[59], p21[59], p22[59], p23[59], p24[59], p25[59], p26[59], p27[59], p28[59], p29[59], p30[59], p31[59], data,data_unq,clk, count59);
 count_mul_v2 x70(p0[60], p1[60], p2[60], p3[60], p4[60], p5[60], p6[60], p7[60], p8[60], p9[60], p10[60], p11[60], p12[60], p13[60], p14[60], p15[60], p16[60], p17[60], p18[60], p19[60], p20[60], p21[60], p22[60], p23[60], p24[60], p25[60], p26[60], p27[60], p28[60], p29[60], p30[60], p31[60], data,data_unq,clk, count60);
 count_mul_v2 x71(p0[61], p1[61], p2[61], p3[61], p4[61], p5[61], p6[61], p7[61], p8[61], p9[61], p10[61], p11[61], p12[61], p13[61], p14[61], p15[61], p16[61], p17[61], p18[61], p19[61], p20[61], p21[61], p22[61], p23[61], p24[61], p25[61], p26[61], p27[61], p28[61], p29[61], p30[61], p31[61], data,data_unq,clk, count61);
 count_mul_v2 x72(p0[62], p1[62], p2[62], p3[62], p4[62], p5[62], p6[62], p7[62], p8[62], p9[62], p10[62], p11[62], p12[62], p13[62], p14[62], p15[62], p16[62], p17[62], p18[62], p19[62], p20[62], p21[62], p22[62], p23[62], p24[62], p25[62], p26[62], p27[62], p28[62], p29[62], p30[62], p31[62], data,data_unq,clk, count62);
 count_mul_v2 x73(p0[63], p1[63], p2[63], p3[63], p4[63], p5[63], p6[63], p7[63], p8[63], p9[63], p10[63], p11[63], p12[63], p13[63], p14[63], p15[63], p16[63], p17[63], p18[63], p19[63], p20[63], p21[63], p22[63], p23[63], p24[63], p25[63], p26[63], p27[63], p28[63], p29[63], p30[63], p31[63], data,data_unq,clk, count63);
 
 
 
 /*
 #include <stdio.h>
 
 int main() {
     // Write C code here
     for (int i = 0; i<64; i++){
     printf("count_ones_new x%d(p0[%d], p1[%d], p2[%d], p3[%d], p4[%d], p5[%d], p6[%d], p7[%d], p8[%d], p9[%d], p10[%d], p11[%d], p12[%d], p13[%d], p14[%d], p15[%d], p16[%d], p17[%d], p18[%d], p19[%d], p20[%d], p21[%d], p22[%d], p23[%d], p24[%d], p25[%d], p26[%d], p27[%d], p28[%d], p29[%d], p30[%d], p31[%d], data,data_unq,clk, count%d); \n\r",10+i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i,i);
     }
 
     return 0;
 }

 
 */
 
 assign pps0 = {count63[0], count62[0], count61[0], count60[0], count59[0], count58[0], count57[0], count56[0], count55[0], count54[0], count53[0], count52[0], count51[0], count50[0], count49[0], count48[0], count47[0], count46[0], count45[0], count44[0], count43[0], count42[0], count41[0], count40[0], count39[0], count38[0], count37[0], count36[0], count35[0], count34[0], count33[0], count32[0], count31[0], count30[0], count29[0], count28[0], count27[0], count26[0], count25[0], count24[0], count23[0], count22[0], count21[0], count20[0], count19[0], count18[0], count17[0], count16[0], count15[0], count14[0], count13[0], count12[0], count11[0], count10[0], count9[0], count8[0], count7[0], count6[0], count5[0], count4[0], count3[0], count2[0], count1[0], count0[0]};
 assign pps1 = {count63[1], count62[1], count61[1], count60[1], count59[1], count58[1], count57[1], count56[1], count55[1], count54[1], count53[1], count52[1], count51[1], count50[1], count49[1], count48[1], count47[1], count46[1], count45[1], count44[1], count43[1], count42[1], count41[1], count40[1], count39[1], count38[1], count37[1], count36[1], count35[1], count34[1], count33[1], count32[1], count31[1], count30[1], count29[1], count28[1], count27[1], count26[1], count25[1], count24[1], count23[1], count22[1], count21[1], count20[1], count19[1], count18[1], count17[1], count16[1], count15[1], count14[1], count13[1], count12[1], count11[1], count10[1], count9[1], count8[1], count7[1], count6[1], count5[1], count4[1], count3[1], count2[1], count1[1], count0[1], 1'b0}; // sum = {sum,count0[0]}
 assign pps2 = {count63[2], count62[2], count61[2], count60[2], count59[2], count58[2], count57[2], count56[2], count55[2], count54[2], count53[2], count52[2], count51[2], count50[2], count49[2], count48[2], count47[2], count46[2], count45[2], count44[2], count43[2], count42[2], count41[2], count40[2], count39[2], count38[2], count37[2], count36[2], count35[2], count34[2], count33[2], count32[2], count31[2], count30[2], count29[2], count28[2], count27[2], count26[2], count25[2], count24[2], count23[2], count22[2], count21[2], count20[2], count19[2], count18[2], count17[2], count16[2], count15[2], count14[2], count13[2], count12[2], count11[2], count10[2], count9[2], count8[2], count7[2], count6[2], count5[2], count4[2], count3[2], count2[2], count1[2], count0[2], 1'b0, 1'b0};
 assign pps3 = {count63[3], count62[3], count61[3], count60[3], count59[3], count58[3], count57[3], count56[3], count55[3], count54[3], count53[3], count52[3], count51[3], count50[3], count49[3], count48[3], count47[3], count46[3], count45[3], count44[3], count43[3], count42[3], count41[3], count40[3], count39[3], count38[3], count37[3], count36[3], count35[3], count34[3], count33[3], count32[3], count31[3], count30[3], count29[3], count28[3], count27[3], count26[3], count25[3], count24[3], count23[3], count22[3], count21[3], count20[3], count19[3], count18[3], count17[3], count16[3], count15[3], count14[3], count13[3], count12[3], count11[3], count10[3], count9[3], count8[3], count7[3], count6[3], count5[3], count4[3], count3[3], count2[3], count1[3], count0[3], 1'b0, 1'b0, 1'b0};// sum = {sum,count0[2],1'b0,1'b0}
 assign pps4=  {count63[4], count62[4], count61[4], count60[4], count59[4], count58[4], count57[4], count56[4], count55[4], count54[4], count53[4], count52[4], count51[4], count50[4], count49[4], count48[4], count47[4], count46[4], count45[4], count44[4], count43[4], count42[4], count41[4], count40[4], count39[4], count38[4], count37[4], count36[4], count35[4], count34[4], count33[4], count32[4], count31[4], count30[4], count29[4], count28[4], count27[4], count26[4], count25[4], count24[4], count23[4], count22[4], count21[4], count20[4], count19[4], count18[4], count17[4], count16[4], count15[4], count14[4], count13[4], count12[4], count11[4], count10[4], count9[4], count8[4], count7[4], count6[4], count5[4], count4[4], count3[4], count2[4], count1[4], count0[4], 1'b0, 1'b0, 1'b0, 1'b0};// sum = {sum,count0[4],1'b0,1'b0,1'b0,1'b0}
 assign pps5 = {count63[5], count62[5], count61[5], count60[5], count59[5], count58[5], count57[5], count56[5], count55[5], count54[5], count53[5], count52[5], count51[5], count50[5], count49[5], count48[5], count47[5], count46[5], count45[5], count44[5], count43[5], count42[5], count41[5], count40[5], count39[5], count38[5], count37[5], count36[5], count35[5], count34[5], count33[5], count32[5], count31[5], count30[5], count29[5], count28[5], count27[5], count26[5], count25[5], count24[5], count23[5], count22[5], count21[5], count20[5], count19[5], count18[5], count17[5], count16[5], count15[5], count14[5], count13[5], count12[5], count11[5], count10[5], count9[5], count8[5], count7[5], count6[5], count5[5], count4[5], count3[5], count2[5], count1[5], count0[5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}; //69 bit width
 /////// OBJECTIVE is : ppso+pps1+pps2+pps3+pps4+pps5
 assign actualsum_pps = pps0+pps1+pps2+pps3+pps4+pps5;
 
adder_64bit_re mod_ad64_0(clk,rst,1'b1,{1'b0,pps0[63:1]},pps1[64:1],64'b0,data,data_unq,sum_pps01,actual_sum01,final_flag01); // sum = {sum,count0[0]}
adder_64bit_re mod_ad64_1(clk,rst,1'b1,{1'b0,pps2[65:3]},pps3[66:3],64'b0,data,data_unq,sum_pps23,actual_sum23,final_flag23);// sum = {sum,count0[2],1'b0,1'b0}
adder_64bit_re mod_ad64_2(clk,rst,1'b1,{1'b0,pps4[67:5]},pps5[68:5],64'b0,data,data_unq,sum_pps45,actual_sum45,final_flag45);// sum = {sum,count0[4],1'b0,1'b0,1'b0,1'b0}

adder_68bit_re mod_ad68_0(clk,rst,1'b1,{ 1'b0, 1'b0,sum_pps01, count0[0]},{sum_pps23, count0[2], 1'b0, 1'b0},68'b0,data,data_unq,sum_pps0123,actual_sum0123,final_flag0123);// sum = {sum,count0[4],1'b0,1'b0,1'b0,1'b0}
adder_72bit_re mod_ad72_0(clk,rst,1'b1,{1'b0,1'b0,sum_pps45, count0[4], 1'b0, 1'b0, 1'b0, 1'b0},{1'b0,1'b0,1'b0,sum_pps0123},72'b0,data,data_unq,sum_pps012345,actual_sum012345,final_flag012345);// sum = {sum,count0[4],1'b0,1'b0,1'b0,1'b0}



//adder_68bit_re mod_ad72_0(clk,rst,1'b1,sum_pps45[63:0],sum_pps0123[63:0],72'b0,data,data_unq,sum_pps012345,actual_sum012345,final_flag012345);// sum = {sum,count0[4],1'b0,1'b0,1'b0,1'b0}



assign sum = sum_pps012345;



assign actualsum_pps01_23_45 = 
    {sum_pps01, count0[0]} + //65bit
    {sum_pps23, count0[2], 1'b0, 1'b0} +  //68bit
    {sum_pps45, count0[4], 1'b0, 1'b0, 1'b0, 1'b0}; //72bit

//assign sum = {actualsum_pps01_23_45,sum_pps01[0],count0[0]};







 /*
 
 assign ppk0 = { 
     sum16_ppk0[4:0], 
     sum15_ppk0[3:0], 
     sum14_ppk0[3:0], 
     sum13_ppk0[3:0], 
     sum12_ppk0[3:0], 
     sum11_ppk0[3:0], 
     sum10_ppk0[3:0], 
     sum9_ppk0[3:0], 
     sum8_ppk0[3:0], 
     sum7_ppk0[3:0], 
     sum6_ppk0[3:0], 
     sum5_ppk0[3:0], 
     sum4_ppk0[3:0], 
     sum3_ppk0[3:0], 
     sum2_ppk0[3:0], 
     sum1_ppk0[3:0], 
     sum0_ppk0[3:0]
 };
 */
endmodule



module multiplier(
input logic [31:0] A,B,
input logic  clk,
output logic [63:0] out
    );
    logic data_flag;
    logic [1:0] and_op [7:0]; // CAM cell 
    logic addr[1024];
    logic loop_0 ,loop_1 ,loop_2 ,loop_3 ,loop_4 ,loop_5 ,loop_6 ,loop_7 ,loop_8 ,loop_9 ,loop_10 ,loop_11 ,loop_12 ,loop_13 ,loop_14 ,loop_15 ,loop_16 ,loop_17 ,loop_18 ,loop_19 ,loop_20 ,loop_21 ,loop_22 ,loop_23 ,loop_24 ,loop_25 ,loop_26 ,loop_27 ,loop_28 ,loop_29 ,loop_30 ,loop_31 ,loop_32 ,loop_33 ,loop_34 ,loop_35 ,loop_36 ,loop_37 ,loop_38 ,loop_39 ,loop_40 ,loop_41 ,loop_42 ,loop_43 ,loop_44 ,loop_45 ,loop_46 ,loop_47 ,loop_48 ,loop_49 ,loop_50 ,loop_51 ,loop_52 ,loop_53 ,loop_54 ,loop_55 ,loop_56 ,loop_57 ,loop_58 ,loop_59 ,loop_60 ,loop_61 ,loop_62 ,loop_63 ,loop_64 ,loop_65 ,loop_66 ,loop_67 ,loop_68 ,loop_69 ,loop_70 ,loop_71 ,loop_72 ,loop_73 ,loop_74 ,loop_75 ,loop_76 ,loop_77 ,loop_78 ,loop_79 ,loop_80 ,loop_81 ,loop_82 ,loop_83 ,loop_84 ,loop_85 ,loop_86 ,loop_87 ,loop_88 ,loop_89 ,loop_90 ,loop_91 ,loop_92 ,loop_93 ,loop_94 ,loop_95 ,loop_96 ,loop_97 ,loop_98 ,loop_99 ,loop_100 ,loop_101 ,loop_102 ,loop_103 ,loop_104 ,loop_105 ,loop_106 ,loop_107 ,loop_108 ,loop_109 ,loop_110 ,loop_111 ,loop_112 ,loop_113 ,loop_114 ,loop_115 ,loop_116 ,loop_117 ,loop_118 ,loop_119 ,loop_120 ,loop_121 ,loop_122 ,loop_123 ,loop_124 ,loop_125 ,loop_126 ,loop_127 ,loop_128 ,loop_129 ,loop_130 ,loop_131 ,loop_132 ,loop_133 ,loop_134 ,loop_135 ,loop_136 ,loop_137 ,loop_138 ,loop_139 ,loop_140 ,loop_141 ,loop_142 ,loop_143 ,loop_144 ,loop_145 ,loop_146 ,loop_147 ,loop_148 ,loop_149 ,loop_150 ,loop_151 ,loop_152 ,loop_153 ,loop_154 ,loop_155 ,loop_156 ,loop_157 ,loop_158 ,loop_159 ,loop_160 ,loop_161 ,loop_162 ,loop_163 ,loop_164 ,loop_165 ,loop_166 ,loop_167 ,loop_168 ,loop_169 ,loop_170 ,loop_171 ,loop_172 ,loop_173 ,loop_174 ,loop_175 ,loop_176 ,loop_177 ,loop_178 ,loop_179 ,loop_180 ,loop_181 ,loop_182 ,loop_183 ,loop_184 ,loop_185 ,loop_186 ,loop_187 ,loop_188 ,loop_189 ,loop_190 ,loop_191 ,loop_192 ,loop_193 ,loop_194 ,loop_195 ,loop_196 ,loop_197 ,loop_198 ,loop_199 ,loop_200 ,loop_201 ,loop_202 ,loop_203 ,loop_204 ,loop_205 ,loop_206 ,loop_207 ,loop_208 ,loop_209 ,loop_210 ,loop_211 ,loop_212 ,loop_213 ,loop_214 ,loop_215 ,loop_216 ,loop_217 ,loop_218 ,loop_219 ,loop_220 ,loop_221 ,loop_222 ,loop_223 ,loop_224 ,loop_225 ,loop_226 ,loop_227 ,loop_228 ,loop_229 ,loop_230 ,loop_231 ,loop_232 ,loop_233 ,loop_234 ,loop_235 ,loop_236 ,loop_237 ,loop_238 ,loop_239 ,loop_240 ,loop_241 ,loop_242 ,loop_243 ,loop_244 ,loop_245 ,loop_246 ,loop_247 ,loop_248 ,loop_249 ,loop_250 ,loop_251 ,loop_252 ,loop_253 ,loop_254 ,loop_255 ,loop_256 ,loop_257 ,loop_258 ,loop_259 ,loop_260 ,loop_261 ,loop_262 ,loop_263 ,loop_264 ,loop_265 ,loop_266 ,loop_267 ,loop_268 ,loop_269 ,loop_270 ,loop_271 ,loop_272 ,loop_273 ,loop_274 ,loop_275 ,loop_276 ,loop_277 ,loop_278 ,loop_279 ,loop_280 ,loop_281 ,loop_282 ,loop_283 ,loop_284 ,loop_285 ,loop_286 ,loop_287 ,loop_288 ,loop_289 ,loop_290 ,loop_291 ,loop_292 ,loop_293 ,loop_294 ,loop_295 ,loop_296 ,loop_297 ,loop_298 ,loop_299 ,loop_300 ,loop_301 ,loop_302 ,loop_303 ,loop_304 ,loop_305 ,loop_306 ,loop_307 ,loop_308 ,loop_309 ,loop_310 ,loop_311 ,loop_312 ,loop_313 ,loop_314 ,loop_315 ,loop_316 ,loop_317 ,loop_318 ,loop_319 ,loop_320 ,loop_321 ,loop_322 ,loop_323 ,loop_324 ,loop_325 ,loop_326 ,loop_327 ,loop_328 ,loop_329 ,loop_330 ,loop_331 ,loop_332 ,loop_333 ,loop_334 ,loop_335 ,loop_336 ,loop_337 ,loop_338 ,loop_339 ,loop_340 ,loop_341 ,loop_342 ,loop_343 ,loop_344 ,loop_345 ,loop_346 ,loop_347 ,loop_348 ,loop_349 ,loop_350 ,loop_351 ,loop_352 ,loop_353 ,loop_354 ,loop_355 ,loop_356 ,loop_357 ,loop_358 ,loop_359 ,loop_360 ,loop_361 ,loop_362 ,loop_363 ,loop_364 ,loop_365 ,loop_366 ,loop_367 ,loop_368 ,loop_369 ,loop_370 ,loop_371 ,loop_372 ,loop_373 ,loop_374 ,loop_375 ,loop_376 ,loop_377 ,loop_378 ,loop_379 ,loop_380 ,loop_381 ,loop_382 ,loop_383 ,loop_384 ,loop_385 ,loop_386 ,loop_387 ,loop_388 ,loop_389 ,loop_390 ,loop_391 ,loop_392 ,loop_393 ,loop_394 ,loop_395 ,loop_396 ,loop_397 ,loop_398 ,loop_399 ,loop_400 ,loop_401 ,loop_402 ,loop_403 ,loop_404 ,loop_405 ,loop_406 ,loop_407 ,loop_408 ,loop_409 ,loop_410 ,loop_411 ,loop_412 ,loop_413 ,loop_414 ,loop_415 ,loop_416 ,loop_417 ,loop_418 ,loop_419 ,loop_420 ,loop_421 ,loop_422 ,loop_423 ,loop_424 ,loop_425 ,loop_426 ,loop_427 ,loop_428 ,loop_429 ,loop_430 ,loop_431 ,loop_432 ,loop_433 ,loop_434 ,loop_435 ,loop_436 ,loop_437 ,loop_438 ,loop_439 ,loop_440 ,loop_441 ,loop_442 ,loop_443 ,loop_444 ,loop_445 ,loop_446 ,loop_447 ,loop_448 ,loop_449 ,loop_450 ,loop_451 ,loop_452 ,loop_453 ,loop_454 ,loop_455 ,loop_456 ,loop_457 ,loop_458 ,loop_459 ,loop_460 ,loop_461 ,loop_462 ,loop_463 ,loop_464 ,loop_465 ,loop_466 ,loop_467 ,loop_468 ,loop_469 ,loop_470 ,loop_471 ,loop_472 ,loop_473 ,loop_474 ,loop_475 ,loop_476 ,loop_477 ,loop_478 ,loop_479 ,loop_480 ,loop_481 ,loop_482 ,loop_483 ,loop_484 ,loop_485 ,loop_486 ,loop_487 ,loop_488 ,loop_489 ,loop_490 ,loop_491 ,loop_492 ,loop_493 ,loop_494 ,loop_495 ,loop_496 ,loop_497 ,loop_498 ,loop_499 ,loop_500 ,loop_501 ,loop_502 ,loop_503 ,loop_504 ,loop_505 ,loop_506 ,loop_507 ,loop_508 ,loop_509 ,loop_510 ,loop_511 ,loop_512 ,loop_513 ,loop_514 ,loop_515 ,loop_516 ,loop_517 ,loop_518 ,loop_519 ,loop_520 ,loop_521 ,loop_522 ,loop_523 ,loop_524 ,loop_525 ,loop_526 ,loop_527 ,loop_528 ,loop_529 ,loop_530 ,loop_531 ,loop_532 ,loop_533 ,loop_534 ,loop_535 ,loop_536 ,loop_537 ,loop_538 ,loop_539 ,loop_540 ,loop_541 ,loop_542 ,loop_543 ,loop_544 ,loop_545 ,loop_546 ,loop_547 ,loop_548 ,loop_549 ,loop_550 ,loop_551 ,loop_552 ,loop_553 ,loop_554 ,loop_555 ,loop_556 ,loop_557 ,loop_558 ,loop_559 ,loop_560 ,loop_561 ,loop_562 ,loop_563 ,loop_564 ,loop_565 ,loop_566 ,loop_567 ,loop_568 ,loop_569 ,loop_570 ,loop_571 ,loop_572 ,loop_573 ,loop_574 ,loop_575 ,loop_576 ,loop_577 ,loop_578 ,loop_579 ,loop_580 ,loop_581 ,loop_582 ,loop_583 ,loop_584 ,loop_585 ,loop_586 ,loop_587 ,loop_588 ,loop_589 ,loop_590 ,loop_591 ,loop_592 ,loop_593 ,loop_594 ,loop_595 ,loop_596 ,loop_597 ,loop_598 ,loop_599 ,loop_600 ,loop_601 ,loop_602 ,loop_603 ,loop_604 ,loop_605 ,loop_606 ,loop_607 ,loop_608 ,loop_609 ,loop_610 ,loop_611 ,loop_612 ,loop_613 ,loop_614 ,loop_615 ,loop_616 ,loop_617 ,loop_618 ,loop_619 ,loop_620 ,loop_621 ,loop_622 ,loop_623 ,loop_624 ,loop_625 ,loop_626 ,loop_627 ,loop_628 ,loop_629 ,loop_630 ,loop_631 ,loop_632 ,loop_633 ,loop_634 ,loop_635 ,loop_636 ,loop_637 ,loop_638 ,loop_639 ,loop_640 ,loop_641 ,loop_642 ,loop_643 ,loop_644 ,loop_645 ,loop_646 ,loop_647 ,loop_648 ,loop_649 ,loop_650 ,loop_651 ,loop_652 ,loop_653 ,loop_654 ,loop_655 ,loop_656 ,loop_657 ,loop_658 ,loop_659 ,loop_660 ,loop_661 ,loop_662 ,loop_663 ,loop_664 ,loop_665 ,loop_666 ,loop_667 ,loop_668 ,loop_669 ,loop_670 ,loop_671 ,loop_672 ,loop_673 ,loop_674 ,loop_675 ,loop_676 ,loop_677 ,loop_678 ,loop_679 ,loop_680 ,loop_681 ,loop_682 ,loop_683 ,loop_684 ,loop_685 ,loop_686 ,loop_687 ,loop_688 ,loop_689 ,loop_690 ,loop_691 ,loop_692 ,loop_693 ,loop_694 ,loop_695 ,loop_696 ,loop_697 ,loop_698 ,loop_699 ,loop_700 ,loop_701 ,loop_702 ,loop_703 ,loop_704 ,loop_705 ,loop_706 ,loop_707 ,loop_708 ,loop_709 ,loop_710 ,loop_711 ,loop_712 ,loop_713 ,loop_714 ,loop_715 ,loop_716 ,loop_717 ,loop_718 ,loop_719 ,loop_720 ,loop_721 ,loop_722 ,loop_723 ,loop_724 ,loop_725 ,loop_726 ,loop_727 ,loop_728 ,loop_729 ,loop_730 ,loop_731 ,loop_732 ,loop_733 ,loop_734 ,loop_735 ,loop_736 ,loop_737 ,loop_738 ,loop_739 ,loop_740 ,loop_741 ,loop_742 ,loop_743 ,loop_744 ,loop_745 ,loop_746 ,loop_747 ,loop_748 ,loop_749 ,loop_750 ,loop_751 ,loop_752 ,loop_753 ,loop_754 ,loop_755 ,loop_756 ,loop_757 ,loop_758 ,loop_759 ,loop_760 ,loop_761 ,loop_762 ,loop_763 ,loop_764 ,loop_765 ,loop_766 ,loop_767 ,loop_768 ,loop_769 ,loop_770 ,loop_771 ,loop_772 ,loop_773 ,loop_774 ,loop_775 ,loop_776 ,loop_777 ,loop_778 ,loop_779 ,loop_780 ,loop_781 ,loop_782 ,loop_783 ,loop_784 ,loop_785 ,loop_786 ,loop_787 ,loop_788 ,loop_789 ,loop_790 ,loop_791 ,loop_792 ,loop_793 ,loop_794 ,loop_795 ,loop_796 ,loop_797 ,loop_798 ,loop_799 ,loop_800 ,loop_801 ,loop_802 ,loop_803 ,loop_804 ,loop_805 ,loop_806 ,loop_807 ,loop_808 ,loop_809 ,loop_810 ,loop_811 ,loop_812 ,loop_813 ,loop_814 ,loop_815 ,loop_816 ,loop_817 ,loop_818 ,loop_819 ,loop_820 ,loop_821 ,loop_822 ,loop_823 ,loop_824 ,loop_825 ,loop_826 ,loop_827 ,loop_828 ,loop_829 ,loop_830 ,loop_831 ,loop_832 ,loop_833 ,loop_834 ,loop_835 ,loop_836 ,loop_837 ,loop_838 ,loop_839 ,loop_840 ,loop_841 ,loop_842 ,loop_843 ,loop_844 ,loop_845 ,loop_846 ,loop_847 ,loop_848 ,loop_849 ,loop_850 ,loop_851 ,loop_852 ,loop_853 ,loop_854 ,loop_855 ,loop_856 ,loop_857 ,loop_858 ,loop_859 ,loop_860 ,loop_861 ,loop_862 ,loop_863 ,loop_864 ,loop_865 ,loop_866 ,loop_867 ,loop_868 ,loop_869 ,loop_870 ,loop_871 ,loop_872 ,loop_873 ,loop_874 ,loop_875 ,loop_876 ,loop_877 ,loop_878 ,loop_879 ,loop_880 ,loop_881 ,loop_882 ,loop_883 ,loop_884 ,loop_885 ,loop_886 ,loop_887 ,loop_888 ,loop_889 ,loop_890 ,loop_891 ,loop_892 ,loop_893 ,loop_894 ,loop_895 ,loop_896 ,loop_897 ,loop_898 ,loop_899 ,loop_900 ,loop_901 ,loop_902 ,loop_903 ,loop_904 ,loop_905 ,loop_906 ,loop_907 ,loop_908 ,loop_909 ,loop_910 ,loop_911 ,loop_912 ,loop_913 ,loop_914 ,loop_915 ,loop_916 ,loop_917 ,loop_918 ,loop_919 ,loop_920 ,loop_921 ,loop_922 ,loop_923 ,loop_924 ,loop_925 ,loop_926 ,loop_927 ,loop_928 ,loop_929 ,loop_930 ,loop_931 ,loop_932 ,loop_933 ,loop_934 ,loop_935 ,loop_936 ,loop_937 ,loop_938 ,loop_939 ,loop_940 ,loop_941 ,loop_942 ,loop_943 ,loop_944 ,loop_945 ,loop_946 ,loop_947 ,loop_948 ,loop_949 ,loop_950 ,loop_951 ,loop_952 ,loop_953 ,loop_954 ,loop_955 ,loop_956 ,loop_957 ,loop_958 ,loop_959 ,loop_960 ,loop_961 ,loop_962 ,loop_963 ,loop_964 ,loop_965 ,loop_966 ,loop_967 ,loop_968 ,loop_969 ,loop_970 ,loop_971 ,loop_972 ,loop_973 ,loop_974 ,loop_975 ,loop_976 ,loop_977 ,loop_978 ,loop_979 ,loop_980 ,loop_981 ,loop_982 ,loop_983 ,loop_984 ,loop_985 ,loop_986 ,loop_987 ,loop_988 ,loop_989 ,loop_990 ,loop_991 ,loop_992 ,loop_993 ,loop_994 ,loop_995 ,loop_996 ,loop_997 ,loop_998 ,loop_999 ,loop_1000 ,loop_1001 ,loop_1002 ,loop_1003 ,loop_1004 ,loop_1005 ,loop_1006 ,loop_1007 ,loop_1008 ,loop_1009 ,loop_1010 ,loop_1011 ,loop_1012 ,loop_1013 ,loop_1014 ,loop_1015 ,loop_1016 ,loop_1017 ,loop_1018 ,loop_1019 ,loop_1020 ,loop_1021 ,loop_1022 ,loop_1023;


    logic match_flag_0 ,match_flag_1 ,match_flag_2 ,match_flag_3 ,match_flag_4 ,match_flag_5 ,match_flag_6 ,match_flag_7 
,match_flag_8 ,match_flag_9 ,match_flag_10 ,match_flag_11 ,match_flag_12 ,match_flag_13 ,match_flag_14 ,match_flag_15 
,match_flag_16 ,match_flag_17 ,match_flag_18 ,match_flag_19 ,match_flag_20 ,match_flag_21 ,match_flag_22 ,match_flag_23 
,match_flag_24 ,match_flag_25 ,match_flag_26 ,match_flag_27 ,match_flag_28 ,match_flag_29 ,match_flag_30 ,match_flag_31 
,match_flag_32 ,match_flag_33 ,match_flag_34 ,match_flag_35 ,match_flag_36 ,match_flag_37 ,match_flag_38 ,match_flag_39 
,match_flag_40 ,match_flag_41 ,match_flag_42 ,match_flag_43 ,match_flag_44 ,match_flag_45 ,match_flag_46 ,match_flag_47 
,match_flag_48 ,match_flag_49 ,match_flag_50 ,match_flag_51 ,match_flag_52 ,match_flag_53 ,match_flag_54 ,match_flag_55 
,match_flag_56 ,match_flag_57 ,match_flag_58 ,match_flag_59 ,match_flag_60 ,match_flag_61 ,match_flag_62 ,match_flag_63 
,match_flag_64 ,match_flag_65 ,match_flag_66 ,match_flag_67 ,match_flag_68 ,match_flag_69 ,match_flag_70 ,match_flag_71 
,match_flag_72 ,match_flag_73 ,match_flag_74 ,match_flag_75 ,match_flag_76 ,match_flag_77 ,match_flag_78 ,match_flag_79 
,match_flag_80 ,match_flag_81 ,match_flag_82 ,match_flag_83 ,match_flag_84 ,match_flag_85 ,match_flag_86 ,match_flag_87 
,match_flag_88 ,match_flag_89 ,match_flag_90 ,match_flag_91 ,match_flag_92 ,match_flag_93 ,match_flag_94 ,match_flag_95 
,match_flag_96 ,match_flag_97 ,match_flag_98 ,match_flag_99 ,match_flag_100 ,match_flag_101 ,match_flag_102 ,match_flag_103 
,match_flag_104 ,match_flag_105 ,match_flag_106 ,match_flag_107 ,match_flag_108 ,match_flag_109 ,match_flag_110 ,match_flag_111 
,match_flag_112 ,match_flag_113 ,match_flag_114 ,match_flag_115 ,match_flag_116 ,match_flag_117 ,match_flag_118 ,match_flag_119 
,match_flag_120 ,match_flag_121 ,match_flag_122 ,match_flag_123 ,match_flag_124 ,match_flag_125 ,match_flag_126 ,match_flag_127 
,match_flag_128 ,match_flag_129 ,match_flag_130 ,match_flag_131 ,match_flag_132 ,match_flag_133 ,match_flag_134 ,match_flag_135 
,match_flag_136 ,match_flag_137 ,match_flag_138 ,match_flag_139 ,match_flag_140 ,match_flag_141 ,match_flag_142 ,match_flag_143
 ,match_flag_144 ,match_flag_145 ,match_flag_146 ,match_flag_147 ,match_flag_148 ,match_flag_149 ,match_flag_150 ,match_flag_151
 ,match_flag_152 ,match_flag_153 ,match_flag_154 ,match_flag_155 ,match_flag_156 ,match_flag_157 ,match_flag_158 ,match_flag_159 ,match_flag_160 ,match_flag_161 ,match_flag_162 ,match_flag_163 ,match_flag_164 ,match_flag_165 ,match_flag_166 ,match_flag_167 ,match_flag_168 ,match_flag_169 ,match_flag_170 ,match_flag_171 ,match_flag_172 ,match_flag_173 ,match_flag_174 ,match_flag_175 ,match_flag_176 ,match_flag_177 ,match_flag_178 ,match_flag_179 ,match_flag_180 ,match_flag_181 ,match_flag_182 ,match_flag_183 ,match_flag_184 ,match_flag_185 ,match_flag_186 ,match_flag_187 ,match_flag_188 ,match_flag_189 ,match_flag_190 ,match_flag_191 ,match_flag_192 ,match_flag_193 ,match_flag_194 ,match_flag_195 ,match_flag_196 ,match_flag_197 ,match_flag_198 ,match_flag_199 ,match_flag_200 ,match_flag_201 ,match_flag_202 ,match_flag_203 ,match_flag_204 ,match_flag_205 ,match_flag_206 ,match_flag_207 ,match_flag_208 ,match_flag_209 ,match_flag_210 ,match_flag_211 ,match_flag_212 ,match_flag_213 ,match_flag_214 ,match_flag_215 ,match_flag_216 ,match_flag_217 ,match_flag_218 ,match_flag_219 ,match_flag_220 ,match_flag_221 ,match_flag_222 ,match_flag_223 ,match_flag_224 ,match_flag_225 ,match_flag_226 ,match_flag_227 ,match_flag_228 ,match_flag_229 ,match_flag_230 ,match_flag_231 ,match_flag_232 ,match_flag_233 ,match_flag_234 ,match_flag_235 ,match_flag_236 ,match_flag_237 ,match_flag_238 ,match_flag_239 ,match_flag_240 ,match_flag_241 ,match_flag_242 ,match_flag_243 ,match_flag_244 ,match_flag_245 ,match_flag_246 ,match_flag_247 ,match_flag_248 ,match_flag_249 ,match_flag_250 ,match_flag_251 ,match_flag_252 ,match_flag_253 ,match_flag_254 ,match_flag_255 ,match_flag_256 ,match_flag_257 ,match_flag_258 ,match_flag_259 ,match_flag_260 ,match_flag_261 ,match_flag_262 ,match_flag_263 ,match_flag_264 ,match_flag_265 ,match_flag_266 ,match_flag_267 ,match_flag_268 ,match_flag_269 ,match_flag_270 ,match_flag_271 ,match_flag_272 ,match_flag_273 ,match_flag_274 ,match_flag_275 ,match_flag_276 ,match_flag_277 ,match_flag_278 ,match_flag_279 ,match_flag_280 ,match_flag_281 ,match_flag_282 ,match_flag_283 ,match_flag_284 ,match_flag_285 ,match_flag_286 ,match_flag_287 ,match_flag_288 ,match_flag_289 ,match_flag_290 ,match_flag_291 ,match_flag_292 ,match_flag_293 ,match_flag_294 ,match_flag_295 ,match_flag_296 ,match_flag_297 ,match_flag_298 ,match_flag_299 ,match_flag_300 ,match_flag_301 ,match_flag_302 ,match_flag_303 ,match_flag_304 ,match_flag_305 ,match_flag_306 ,match_flag_307 ,match_flag_308 ,match_flag_309 ,match_flag_310 ,match_flag_311 ,match_flag_312 ,match_flag_313 ,match_flag_314 ,match_flag_315 ,match_flag_316 ,match_flag_317 ,match_flag_318 ,match_flag_319 ,match_flag_320 ,match_flag_321 ,match_flag_322 ,match_flag_323 ,match_flag_324 ,match_flag_325 ,match_flag_326 ,match_flag_327 ,match_flag_328 ,match_flag_329 ,match_flag_330 ,match_flag_331 ,match_flag_332 ,match_flag_333 ,match_flag_334 ,match_flag_335 ,match_flag_336 ,match_flag_337 ,match_flag_338 ,match_flag_339 ,match_flag_340 ,match_flag_341 ,match_flag_342 ,match_flag_343 ,match_flag_344 ,match_flag_345 ,match_flag_346 ,match_flag_347 ,match_flag_348 ,match_flag_349 ,match_flag_350 ,match_flag_351 ,match_flag_352 ,match_flag_353 ,match_flag_354 ,match_flag_355 ,match_flag_356 ,match_flag_357 ,match_flag_358 ,match_flag_359 ,match_flag_360 ,match_flag_361 ,match_flag_362 ,match_flag_363 ,match_flag_364 ,match_flag_365 ,match_flag_366 ,match_flag_367 ,match_flag_368 ,match_flag_369 ,match_flag_370 ,match_flag_371 ,match_flag_372 ,match_flag_373 ,match_flag_374 ,match_flag_375 ,match_flag_376 ,match_flag_377 ,match_flag_378 ,match_flag_379 ,match_flag_380 ,match_flag_381 ,match_flag_382 ,match_flag_383 ,match_flag_384 ,match_flag_385 ,match_flag_386 ,match_flag_387 ,match_flag_388 ,match_flag_389 ,match_flag_390 ,match_flag_391 ,match_flag_392 ,match_flag_393 ,match_flag_394 ,match_flag_395 ,match_flag_396 ,match_flag_397 ,match_flag_398 ,match_flag_399 ,match_flag_400 ,match_flag_401 ,match_flag_402 ,match_flag_403 ,match_flag_404 ,match_flag_405 ,match_flag_406 ,match_flag_407 ,match_flag_408 ,match_flag_409 ,match_flag_410 ,match_flag_411 ,match_flag_412 ,match_flag_413 ,match_flag_414 ,match_flag_415 ,match_flag_416 ,match_flag_417 ,match_flag_418 ,match_flag_419 ,match_flag_420 ,match_flag_421 ,match_flag_422 ,match_flag_423 ,match_flag_424 ,match_flag_425 ,match_flag_426 ,match_flag_427 ,match_flag_428 ,match_flag_429 ,match_flag_430 ,match_flag_431 ,match_flag_432 ,match_flag_433 ,match_flag_434 ,match_flag_435 ,match_flag_436 ,match_flag_437 ,match_flag_438 ,match_flag_439 ,match_flag_440 ,match_flag_441 ,match_flag_442 ,match_flag_443 ,match_flag_444 ,match_flag_445 ,match_flag_446 ,match_flag_447 ,match_flag_448 ,match_flag_449 ,match_flag_450 ,match_flag_451 ,match_flag_452 ,match_flag_453 ,match_flag_454 ,match_flag_455 ,match_flag_456 ,match_flag_457 ,match_flag_458 ,match_flag_459 ,match_flag_460 ,match_flag_461 ,match_flag_462 ,match_flag_463 ,match_flag_464 ,match_flag_465 ,match_flag_466 ,match_flag_467 ,match_flag_468 ,match_flag_469 ,match_flag_470 ,match_flag_471 ,match_flag_472 ,match_flag_473 ,match_flag_474 ,match_flag_475 ,match_flag_476 ,match_flag_477 ,match_flag_478 ,match_flag_479 ,match_flag_480 ,match_flag_481 ,match_flag_482 ,match_flag_483 ,match_flag_484 ,match_flag_485 ,match_flag_486 ,match_flag_487 ,match_flag_488 ,match_flag_489 ,match_flag_490 ,match_flag_491 ,match_flag_492 ,match_flag_493 ,match_flag_494 ,match_flag_495 ,match_flag_496 ,match_flag_497 ,match_flag_498 ,match_flag_499 ,match_flag_500 ,match_flag_501 ,match_flag_502 ,match_flag_503 ,match_flag_504 ,match_flag_505 ,match_flag_506 ,match_flag_507 ,match_flag_508 ,match_flag_509 ,match_flag_510 ,match_flag_511 ,match_flag_512 ,match_flag_513 ,match_flag_514 ,match_flag_515 ,match_flag_516 ,match_flag_517 ,match_flag_518 ,match_flag_519 ,match_flag_520 ,match_flag_521 ,match_flag_522 ,match_flag_523 ,match_flag_524 ,match_flag_525 ,match_flag_526 ,match_flag_527 ,match_flag_528 ,match_flag_529 ,match_flag_530 ,match_flag_531 ,match_flag_532 ,match_flag_533 ,match_flag_534 ,match_flag_535 ,match_flag_536 ,match_flag_537 ,match_flag_538 ,match_flag_539 ,match_flag_540 ,match_flag_541 ,match_flag_542 ,match_flag_543 ,match_flag_544 ,match_flag_545 ,match_flag_546 ,match_flag_547 ,match_flag_548 ,match_flag_549 ,match_flag_550 ,match_flag_551 ,match_flag_552 ,match_flag_553 ,match_flag_554 ,match_flag_555 ,match_flag_556 ,match_flag_557 ,match_flag_558 ,match_flag_559 ,match_flag_560 ,match_flag_561 ,match_flag_562 ,match_flag_563 ,match_flag_564 ,match_flag_565 ,match_flag_566 ,match_flag_567 ,match_flag_568 ,match_flag_569 ,match_flag_570 ,match_flag_571 ,match_flag_572 ,match_flag_573 ,match_flag_574 ,match_flag_575 ,match_flag_576 ,match_flag_577 ,match_flag_578 ,match_flag_579 ,match_flag_580 ,match_flag_581 ,match_flag_582 ,match_flag_583 ,match_flag_584 ,match_flag_585 ,match_flag_586 ,match_flag_587 ,match_flag_588 ,match_flag_589 ,match_flag_590 ,match_flag_591 ,match_flag_592 ,match_flag_593 ,match_flag_594 ,match_flag_595 ,match_flag_596 ,match_flag_597 ,match_flag_598 ,match_flag_599 ,match_flag_600 ,match_flag_601 ,match_flag_602 ,match_flag_603 ,match_flag_604 ,match_flag_605 ,match_flag_606 ,match_flag_607 ,match_flag_608 ,match_flag_609 ,match_flag_610 ,match_flag_611 ,match_flag_612 ,match_flag_613 ,match_flag_614 ,match_flag_615 ,match_flag_616 ,match_flag_617 ,match_flag_618 ,match_flag_619 ,match_flag_620 ,match_flag_621 ,match_flag_622 ,match_flag_623 ,match_flag_624 ,match_flag_625 ,match_flag_626 ,match_flag_627 ,match_flag_628 ,match_flag_629 ,match_flag_630 ,match_flag_631 ,match_flag_632 ,match_flag_633 ,match_flag_634 ,match_flag_635 ,match_flag_636 ,match_flag_637 ,match_flag_638 ,match_flag_639 ,match_flag_640 ,match_flag_641 ,match_flag_642 ,match_flag_643 ,match_flag_644 ,match_flag_645 ,match_flag_646 ,match_flag_647 ,match_flag_648 ,match_flag_649 ,match_flag_650 ,match_flag_651 ,match_flag_652 ,match_flag_653 ,match_flag_654 ,match_flag_655 ,match_flag_656 ,match_flag_657 ,match_flag_658 ,match_flag_659 ,match_flag_660 ,match_flag_661 ,match_flag_662 ,match_flag_663 ,match_flag_664 ,match_flag_665 ,match_flag_666 ,match_flag_667 ,match_flag_668 ,match_flag_669 ,match_flag_670 ,match_flag_671 ,match_flag_672 ,match_flag_673 ,match_flag_674 ,match_flag_675 ,match_flag_676 ,match_flag_677 ,match_flag_678 ,match_flag_679 ,match_flag_680 ,match_flag_681 ,match_flag_682 ,match_flag_683 ,match_flag_684 ,match_flag_685 ,match_flag_686 ,match_flag_687 ,match_flag_688 ,match_flag_689 ,match_flag_690 ,match_flag_691 ,match_flag_692 ,match_flag_693 ,match_flag_694 ,match_flag_695 ,match_flag_696 ,match_flag_697 ,match_flag_698 ,match_flag_699 ,match_flag_700 ,match_flag_701 ,match_flag_702 ,match_flag_703 ,match_flag_704 ,match_flag_705 ,match_flag_706 ,match_flag_707 ,match_flag_708 ,match_flag_709 ,match_flag_710 ,match_flag_711 ,match_flag_712 ,match_flag_713 ,match_flag_714 ,match_flag_715 ,match_flag_716 ,match_flag_717 ,match_flag_718 ,match_flag_719 ,match_flag_720 ,match_flag_721 ,match_flag_722 ,match_flag_723 ,match_flag_724 ,match_flag_725 ,match_flag_726 ,match_flag_727 ,match_flag_728 ,match_flag_729 ,match_flag_730 ,match_flag_731 ,match_flag_732 ,match_flag_733 ,match_flag_734 ,match_flag_735 ,match_flag_736 ,match_flag_737 ,match_flag_738 ,match_flag_739 ,match_flag_740 ,match_flag_741 ,match_flag_742 ,match_flag_743 ,match_flag_744 ,match_flag_745 ,match_flag_746 ,match_flag_747 ,match_flag_748 ,match_flag_749 ,match_flag_750 ,match_flag_751 ,match_flag_752 ,match_flag_753 ,match_flag_754 ,match_flag_755 ,match_flag_756 ,match_flag_757 ,match_flag_758 ,match_flag_759 ,match_flag_760 ,match_flag_761 ,match_flag_762 ,match_flag_763 ,match_flag_764 ,match_flag_765 ,match_flag_766 ,match_flag_767 ,match_flag_768 ,match_flag_769 ,match_flag_770 ,match_flag_771 ,match_flag_772 ,match_flag_773 ,match_flag_774 ,match_flag_775 ,match_flag_776 ,match_flag_777 ,match_flag_778 ,match_flag_779 ,match_flag_780 ,match_flag_781 ,match_flag_782 ,match_flag_783 ,match_flag_784 ,match_flag_785 ,match_flag_786 ,match_flag_787 ,match_flag_788 ,match_flag_789 ,match_flag_790 ,match_flag_791 ,match_flag_792 ,match_flag_793 ,match_flag_794 ,match_flag_795 ,match_flag_796 ,match_flag_797 ,match_flag_798 ,match_flag_799 ,match_flag_800 ,match_flag_801 ,match_flag_802 ,match_flag_803 ,match_flag_804 ,match_flag_805 ,match_flag_806 ,match_flag_807 ,match_flag_808 ,match_flag_809 ,match_flag_810 ,match_flag_811 ,match_flag_812 ,match_flag_813 ,match_flag_814 ,match_flag_815 ,match_flag_816 ,match_flag_817 ,match_flag_818 ,match_flag_819 ,match_flag_820 ,match_flag_821 ,match_flag_822 ,match_flag_823 ,match_flag_824 ,match_flag_825 ,match_flag_826 ,match_flag_827 ,match_flag_828 ,match_flag_829 ,match_flag_830 ,match_flag_831 ,match_flag_832 ,match_flag_833 ,match_flag_834 ,match_flag_835 ,match_flag_836 ,match_flag_837 ,match_flag_838 ,match_flag_839 ,match_flag_840 ,match_flag_841 ,match_flag_842 ,match_flag_843 ,match_flag_844 ,match_flag_845 ,match_flag_846 ,match_flag_847 ,match_flag_848 ,match_flag_849 ,match_flag_850 ,match_flag_851 ,match_flag_852 ,match_flag_853 ,match_flag_854 ,match_flag_855 ,match_flag_856 ,match_flag_857 ,match_flag_858 ,match_flag_859 ,match_flag_860 ,match_flag_861 ,match_flag_862 ,match_flag_863 ,match_flag_864 ,match_flag_865 ,match_flag_866 ,match_flag_867 ,match_flag_868 ,match_flag_869 ,match_flag_870 ,match_flag_871 ,match_flag_872 ,match_flag_873 ,match_flag_874 ,match_flag_875 ,match_flag_876 ,match_flag_877 ,match_flag_878 ,match_flag_879 ,match_flag_880 ,match_flag_881 ,match_flag_882 ,match_flag_883 ,match_flag_884 ,match_flag_885 ,match_flag_886 ,match_flag_887 ,match_flag_888 ,match_flag_889 ,match_flag_890 ,match_flag_891 ,match_flag_892 ,match_flag_893 ,match_flag_894 ,match_flag_895 ,match_flag_896 ,match_flag_897 ,match_flag_898 ,match_flag_899 ,match_flag_900 ,match_flag_901 ,match_flag_902 ,match_flag_903 ,match_flag_904 ,match_flag_905 ,match_flag_906 ,match_flag_907 ,match_flag_908 ,match_flag_909 ,match_flag_910 ,match_flag_911 ,match_flag_912 ,match_flag_913 ,match_flag_914 ,match_flag_915 ,match_flag_916 ,match_flag_917 ,match_flag_918 ,match_flag_919 ,match_flag_920 ,match_flag_921 ,match_flag_922 ,match_flag_923 ,match_flag_924 ,match_flag_925 ,match_flag_926 ,match_flag_927 ,match_flag_928 ,match_flag_929 ,match_flag_930 ,match_flag_931 ,match_flag_932 ,match_flag_933 ,match_flag_934 ,match_flag_935 ,match_flag_936 ,match_flag_937 ,match_flag_938 ,match_flag_939 ,match_flag_940 ,match_flag_941 ,match_flag_942 ,match_flag_943 ,match_flag_944 ,match_flag_945 ,match_flag_946 ,match_flag_947 ,match_flag_948 ,match_flag_949 ,match_flag_950 ,match_flag_951 ,match_flag_952 ,match_flag_953 ,match_flag_954 ,match_flag_955 ,match_flag_956 ,match_flag_957 ,match_flag_958 ,match_flag_959 ,match_flag_960 ,match_flag_961 ,match_flag_962 ,match_flag_963 ,match_flag_964 ,match_flag_965 ,match_flag_966 ,match_flag_967 ,match_flag_968 ,match_flag_969 ,match_flag_970 ,match_flag_971 ,match_flag_972 ,match_flag_973 ,match_flag_974 ,match_flag_975 ,match_flag_976 ,match_flag_977 ,match_flag_978 ,match_flag_979 ,match_flag_980 ,match_flag_981 ,match_flag_982 ,match_flag_983 ,match_flag_984 ,match_flag_985 ,match_flag_986 ,match_flag_987 ,match_flag_988 ,match_flag_989 ,match_flag_990 ,match_flag_991 ,match_flag_992 ,match_flag_993 ,match_flag_994 ,match_flag_995 ,match_flag_996 ,match_flag_997 ,match_flag_998 ,match_flag_999 ,match_flag_1000 ,match_flag_1001 ,match_flag_1002 ,match_flag_1003 ,match_flag_1004 ,match_flag_1005 ,match_flag_1006 ,match_flag_1007 ,match_flag_1008 ,match_flag_1009 ,match_flag_1010 ,match_flag_1011 ,match_flag_1012 ,match_flag_1013 ,match_flag_1014 ,match_flag_1015 ,match_flag_1016 ,match_flag_1017 ,match_flag_1018 ,match_flag_1019 ,match_flag_1020 ,match_flag_1021 ,match_flag_1022 ,match_flag_1023;

 always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_0 = 1'b0;
        addr[0] = 3'b0;
        for (loop_0 = 0; loop_0 < NUM_CELL; loop_0++) begin
         if ({b[0],a[0]}) == loop_0[1:0]) begin
          match_flag_0 = 1'b1;
          addr[0] = loop_0[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1 = 1'b0;
        addr[1] = 3'b0;
        for (loop_1 = 0; loop_1 < NUM_CELL; loop_1++) begin
         if ({b[1],a[0]}) == loop_1[1:0]) begin
          match_flag_1 = 1'b1;
          addr[1] = loop_1[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_2 = 1'b0;
        addr[2] = 3'b0;
        for (loop_2 = 0; loop_2 < NUM_CELL; loop_2++) begin
         if ({b[2],a[0]}) == loop_2[1:0]) begin
          match_flag_2 = 1'b1;
          addr[2] = loop_2[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_3 = 1'b0;
        addr[3] = 3'b0;
        for (loop_3 = 0; loop_3 < NUM_CELL; loop_3++) begin
         if ({b[3],a[0]}) == loop_3[1:0]) begin
          match_flag_3 = 1'b1;
          addr[3] = loop_3[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_4 = 1'b0;
        addr[4] = 3'b0;
        for (loop_4 = 0; loop_4 < NUM_CELL; loop_4++) begin
         if ({b[4],a[0]}) == loop_4[1:0]) begin
          match_flag_4 = 1'b1;
          addr[4] = loop_4[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_5 = 1'b0;
        addr[5] = 3'b0;
        for (loop_5 = 0; loop_5 < NUM_CELL; loop_5++) begin
         if ({b[5],a[0]}) == loop_5[1:0]) begin
          match_flag_5 = 1'b1;
          addr[5] = loop_5[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_6 = 1'b0;
        addr[6] = 3'b0;
        for (loop_6 = 0; loop_6 < NUM_CELL; loop_6++) begin
         if ({b[6],a[0]}) == loop_6[1:0]) begin
          match_flag_6 = 1'b1;
          addr[6] = loop_6[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_7 = 1'b0;
        addr[7] = 3'b0;
        for (loop_7 = 0; loop_7 < NUM_CELL; loop_7++) begin
         if ({b[7],a[0]}) == loop_7[1:0]) begin
          match_flag_7 = 1'b1;
          addr[7] = loop_7[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_8 = 1'b0;
        addr[8] = 3'b0;
        for (loop_8 = 0; loop_8 < NUM_CELL; loop_8++) begin
         if ({b[8],a[0]}) == loop_8[1:0]) begin
          match_flag_8 = 1'b1;
          addr[8] = loop_8[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_9 = 1'b0;
        addr[9] = 3'b0;
        for (loop_9 = 0; loop_9 < NUM_CELL; loop_9++) begin
         if ({b[9],a[0]}) == loop_9[1:0]) begin
          match_flag_9 = 1'b1;
          addr[9] = loop_9[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_10 = 1'b0;
        addr[10] = 3'b0;
        for (loop_10 = 0; loop_10 < NUM_CELL; loop_10++) begin
         if ({b[10],a[0]}) == loop_10[1:0]) begin
          match_flag_10 = 1'b1;
          addr[10] = loop_10[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_11 = 1'b0;
        addr[11] = 3'b0;
        for (loop_11 = 0; loop_11 < NUM_CELL; loop_11++) begin
         if ({b[11],a[0]}) == loop_11[1:0]) begin
          match_flag_11 = 1'b1;
          addr[11] = loop_11[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_12 = 1'b0;
        addr[12] = 3'b0;
        for (loop_12 = 0; loop_12 < NUM_CELL; loop_12++) begin
         if ({b[12],a[0]}) == loop_12[1:0]) begin
          match_flag_12 = 1'b1;
          addr[12] = loop_12[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_13 = 1'b0;
        addr[13] = 3'b0;
        for (loop_13 = 0; loop_13 < NUM_CELL; loop_13++) begin
         if ({b[13],a[0]}) == loop_13[1:0]) begin
          match_flag_13 = 1'b1;
          addr[13] = loop_13[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_14 = 1'b0;
        addr[14] = 3'b0;
        for (loop_14 = 0; loop_14 < NUM_CELL; loop_14++) begin
         if ({b[14],a[0]}) == loop_14[1:0]) begin
          match_flag_14 = 1'b1;
          addr[14] = loop_14[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_15 = 1'b0;
        addr[15] = 3'b0;
        for (loop_15 = 0; loop_15 < NUM_CELL; loop_15++) begin
         if ({b[15],a[0]}) == loop_15[1:0]) begin
          match_flag_15 = 1'b1;
          addr[15] = loop_15[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_16 = 1'b0;
        addr[16] = 3'b0;
        for (loop_16 = 0; loop_16 < NUM_CELL; loop_16++) begin
         if ({b[16],a[0]}) == loop_16[1:0]) begin
          match_flag_16 = 1'b1;
          addr[16] = loop_16[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_17 = 1'b0;
        addr[17] = 3'b0;
        for (loop_17 = 0; loop_17 < NUM_CELL; loop_17++) begin
         if ({b[17],a[0]}) == loop_17[1:0]) begin
          match_flag_17 = 1'b1;
          addr[17] = loop_17[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_18 = 1'b0;
        addr[18] = 3'b0;
        for (loop_18 = 0; loop_18 < NUM_CELL; loop_18++) begin
         if ({b[18],a[0]}) == loop_18[1:0]) begin
          match_flag_18 = 1'b1;
          addr[18] = loop_18[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_19 = 1'b0;
        addr[19] = 3'b0;
        for (loop_19 = 0; loop_19 < NUM_CELL; loop_19++) begin
         if ({b[19],a[0]}) == loop_19[1:0]) begin
          match_flag_19 = 1'b1;
          addr[19] = loop_19[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_20 = 1'b0;
        addr[20] = 3'b0;
        for (loop_20 = 0; loop_20 < NUM_CELL; loop_20++) begin
         if ({b[20],a[0]}) == loop_20[1:0]) begin
          match_flag_20 = 1'b1;
          addr[20] = loop_20[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_21 = 1'b0;
        addr[21] = 3'b0;
        for (loop_21 = 0; loop_21 < NUM_CELL; loop_21++) begin
         if ({b[21],a[0]}) == loop_21[1:0]) begin
          match_flag_21 = 1'b1;
          addr[21] = loop_21[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_22 = 1'b0;
        addr[22] = 3'b0;
        for (loop_22 = 0; loop_22 < NUM_CELL; loop_22++) begin
         if ({b[22],a[0]}) == loop_22[1:0]) begin
          match_flag_22 = 1'b1;
          addr[22] = loop_22[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_23 = 1'b0;
        addr[23] = 3'b0;
        for (loop_23 = 0; loop_23 < NUM_CELL; loop_23++) begin
         if ({b[23],a[0]}) == loop_23[1:0]) begin
          match_flag_23 = 1'b1;
          addr[23] = loop_23[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_24 = 1'b0;
        addr[24] = 3'b0;
        for (loop_24 = 0; loop_24 < NUM_CELL; loop_24++) begin
         if ({b[24],a[0]}) == loop_24[1:0]) begin
          match_flag_24 = 1'b1;
          addr[24] = loop_24[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_25 = 1'b0;
        addr[25] = 3'b0;
        for (loop_25 = 0; loop_25 < NUM_CELL; loop_25++) begin
         if ({b[25],a[0]}) == loop_25[1:0]) begin
          match_flag_25 = 1'b1;
          addr[25] = loop_25[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_26 = 1'b0;
        addr[26] = 3'b0;
        for (loop_26 = 0; loop_26 < NUM_CELL; loop_26++) begin
         if ({b[26],a[0]}) == loop_26[1:0]) begin
          match_flag_26 = 1'b1;
          addr[26] = loop_26[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_27 = 1'b0;
        addr[27] = 3'b0;
        for (loop_27 = 0; loop_27 < NUM_CELL; loop_27++) begin
         if ({b[27],a[0]}) == loop_27[1:0]) begin
          match_flag_27 = 1'b1;
          addr[27] = loop_27[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_28 = 1'b0;
        addr[28] = 3'b0;
        for (loop_28 = 0; loop_28 < NUM_CELL; loop_28++) begin
         if ({b[28],a[0]}) == loop_28[1:0]) begin
          match_flag_28 = 1'b1;
          addr[28] = loop_28[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_29 = 1'b0;
        addr[29] = 3'b0;
        for (loop_29 = 0; loop_29 < NUM_CELL; loop_29++) begin
         if ({b[29],a[0]}) == loop_29[1:0]) begin
          match_flag_29 = 1'b1;
          addr[29] = loop_29[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_30 = 1'b0;
        addr[30] = 3'b0;
        for (loop_30 = 0; loop_30 < NUM_CELL; loop_30++) begin
         if ({b[30],a[0]}) == loop_30[1:0]) begin
          match_flag_30 = 1'b1;
          addr[30] = loop_30[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_31 = 1'b0;
        addr[31] = 3'b0;
        for (loop_31 = 0; loop_31 < NUM_CELL; loop_31++) begin
         if ({b[31],a[0]}) == loop_31[1:0]) begin
          match_flag_31 = 1'b1;
          addr[31] = loop_31[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_32 = 1'b0;
        addr[32] = 3'b0;
        for (loop_32 = 0; loop_32 < NUM_CELL; loop_32++) begin
         if ({b[0],a[1]}) == loop_32[1:0]) begin
          match_flag_32 = 1'b1;
          addr[32] = loop_32[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_33 = 1'b0;
        addr[33] = 3'b0;
        for (loop_33 = 0; loop_33 < NUM_CELL; loop_33++) begin
         if ({b[1],a[1]}) == loop_33[1:0]) begin
          match_flag_33 = 1'b1;
          addr[33] = loop_33[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_34 = 1'b0;
        addr[34] = 3'b0;
        for (loop_34 = 0; loop_34 < NUM_CELL; loop_34++) begin
         if ({b[2],a[1]}) == loop_34[1:0]) begin
          match_flag_34 = 1'b1;
          addr[34] = loop_34[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_35 = 1'b0;
        addr[35] = 3'b0;
        for (loop_35 = 0; loop_35 < NUM_CELL; loop_35++) begin
         if ({b[3],a[1]}) == loop_35[1:0]) begin
          match_flag_35 = 1'b1;
          addr[35] = loop_35[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_36 = 1'b0;
        addr[36] = 3'b0;
        for (loop_36 = 0; loop_36 < NUM_CELL; loop_36++) begin
         if ({b[4],a[1]}) == loop_36[1:0]) begin
          match_flag_36 = 1'b1;
          addr[36] = loop_36[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_37 = 1'b0;
        addr[37] = 3'b0;
        for (loop_37 = 0; loop_37 < NUM_CELL; loop_37++) begin
         if ({b[5],a[1]}) == loop_37[1:0]) begin
          match_flag_37 = 1'b1;
          addr[37] = loop_37[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_38 = 1'b0;
        addr[38] = 3'b0;
        for (loop_38 = 0; loop_38 < NUM_CELL; loop_38++) begin
         if ({b[6],a[1]}) == loop_38[1:0]) begin
          match_flag_38 = 1'b1;
          addr[38] = loop_38[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_39 = 1'b0;
        addr[39] = 3'b0;
        for (loop_39 = 0; loop_39 < NUM_CELL; loop_39++) begin
         if ({b[7],a[1]}) == loop_39[1:0]) begin
          match_flag_39 = 1'b1;
          addr[39] = loop_39[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_40 = 1'b0;
        addr[40] = 3'b0;
        for (loop_40 = 0; loop_40 < NUM_CELL; loop_40++) begin
         if ({b[8],a[1]}) == loop_40[1:0]) begin
          match_flag_40 = 1'b1;
          addr[40] = loop_40[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_41 = 1'b0;
        addr[41] = 3'b0;
        for (loop_41 = 0; loop_41 < NUM_CELL; loop_41++) begin
         if ({b[9],a[1]}) == loop_41[1:0]) begin
          match_flag_41 = 1'b1;
          addr[41] = loop_41[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_42 = 1'b0;
        addr[42] = 3'b0;
        for (loop_42 = 0; loop_42 < NUM_CELL; loop_42++) begin
         if ({b[10],a[1]}) == loop_42[1:0]) begin
          match_flag_42 = 1'b1;
          addr[42] = loop_42[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_43 = 1'b0;
        addr[43] = 3'b0;
        for (loop_43 = 0; loop_43 < NUM_CELL; loop_43++) begin
         if ({b[11],a[1]}) == loop_43[1:0]) begin
          match_flag_43 = 1'b1;
          addr[43] = loop_43[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_44 = 1'b0;
        addr[44] = 3'b0;
        for (loop_44 = 0; loop_44 < NUM_CELL; loop_44++) begin
         if ({b[12],a[1]}) == loop_44[1:0]) begin
          match_flag_44 = 1'b1;
          addr[44] = loop_44[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_45 = 1'b0;
        addr[45] = 3'b0;
        for (loop_45 = 0; loop_45 < NUM_CELL; loop_45++) begin
         if ({b[13],a[1]}) == loop_45[1:0]) begin
          match_flag_45 = 1'b1;
          addr[45] = loop_45[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_46 = 1'b0;
        addr[46] = 3'b0;
        for (loop_46 = 0; loop_46 < NUM_CELL; loop_46++) begin
         if ({b[14],a[1]}) == loop_46[1:0]) begin
          match_flag_46 = 1'b1;
          addr[46] = loop_46[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_47 = 1'b0;
        addr[47] = 3'b0;
        for (loop_47 = 0; loop_47 < NUM_CELL; loop_47++) begin
         if ({b[15],a[1]}) == loop_47[1:0]) begin
          match_flag_47 = 1'b1;
          addr[47] = loop_47[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_48 = 1'b0;
        addr[48] = 3'b0;
        for (loop_48 = 0; loop_48 < NUM_CELL; loop_48++) begin
         if ({b[16],a[1]}) == loop_48[1:0]) begin
          match_flag_48 = 1'b1;
          addr[48] = loop_48[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_49 = 1'b0;
        addr[49] = 3'b0;
        for (loop_49 = 0; loop_49 < NUM_CELL; loop_49++) begin
         if ({b[17],a[1]}) == loop_49[1:0]) begin
          match_flag_49 = 1'b1;
          addr[49] = loop_49[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_50 = 1'b0;
        addr[50] = 3'b0;
        for (loop_50 = 0; loop_50 < NUM_CELL; loop_50++) begin
         if ({b[18],a[1]}) == loop_50[1:0]) begin
          match_flag_50 = 1'b1;
          addr[50] = loop_50[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_51 = 1'b0;
        addr[51] = 3'b0;
        for (loop_51 = 0; loop_51 < NUM_CELL; loop_51++) begin
         if ({b[19],a[1]}) == loop_51[1:0]) begin
          match_flag_51 = 1'b1;
          addr[51] = loop_51[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_52 = 1'b0;
        addr[52] = 3'b0;
        for (loop_52 = 0; loop_52 < NUM_CELL; loop_52++) begin
         if ({b[20],a[1]}) == loop_52[1:0]) begin
          match_flag_52 = 1'b1;
          addr[52] = loop_52[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_53 = 1'b0;
        addr[53] = 3'b0;
        for (loop_53 = 0; loop_53 < NUM_CELL; loop_53++) begin
         if ({b[21],a[1]}) == loop_53[1:0]) begin
          match_flag_53 = 1'b1;
          addr[53] = loop_53[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_54 = 1'b0;
        addr[54] = 3'b0;
        for (loop_54 = 0; loop_54 < NUM_CELL; loop_54++) begin
         if ({b[22],a[1]}) == loop_54[1:0]) begin
          match_flag_54 = 1'b1;
          addr[54] = loop_54[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_55 = 1'b0;
        addr[55] = 3'b0;
        for (loop_55 = 0; loop_55 < NUM_CELL; loop_55++) begin
         if ({b[23],a[1]}) == loop_55[1:0]) begin
          match_flag_55 = 1'b1;
          addr[55] = loop_55[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_56 = 1'b0;
        addr[56] = 3'b0;
        for (loop_56 = 0; loop_56 < NUM_CELL; loop_56++) begin
         if ({b[24],a[1]}) == loop_56[1:0]) begin
          match_flag_56 = 1'b1;
          addr[56] = loop_56[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_57 = 1'b0;
        addr[57] = 3'b0;
        for (loop_57 = 0; loop_57 < NUM_CELL; loop_57++) begin
         if ({b[25],a[1]}) == loop_57[1:0]) begin
          match_flag_57 = 1'b1;
          addr[57] = loop_57[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_58 = 1'b0;
        addr[58] = 3'b0;
        for (loop_58 = 0; loop_58 < NUM_CELL; loop_58++) begin
         if ({b[26],a[1]}) == loop_58[1:0]) begin
          match_flag_58 = 1'b1;
          addr[58] = loop_58[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_59 = 1'b0;
        addr[59] = 3'b0;
        for (loop_59 = 0; loop_59 < NUM_CELL; loop_59++) begin
         if ({b[27],a[1]}) == loop_59[1:0]) begin
          match_flag_59 = 1'b1;
          addr[59] = loop_59[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_60 = 1'b0;
        addr[60] = 3'b0;
        for (loop_60 = 0; loop_60 < NUM_CELL; loop_60++) begin
         if ({b[28],a[1]}) == loop_60[1:0]) begin
          match_flag_60 = 1'b1;
          addr[60] = loop_60[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_61 = 1'b0;
        addr[61] = 3'b0;
        for (loop_61 = 0; loop_61 < NUM_CELL; loop_61++) begin
         if ({b[29],a[1]}) == loop_61[1:0]) begin
          match_flag_61 = 1'b1;
          addr[61] = loop_61[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_62 = 1'b0;
        addr[62] = 3'b0;
        for (loop_62 = 0; loop_62 < NUM_CELL; loop_62++) begin
         if ({b[30],a[1]}) == loop_62[1:0]) begin
          match_flag_62 = 1'b1;
          addr[62] = loop_62[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_63 = 1'b0;
        addr[63] = 3'b0;
        for (loop_63 = 0; loop_63 < NUM_CELL; loop_63++) begin
         if ({b[31],a[1]}) == loop_63[1:0]) begin
          match_flag_63 = 1'b1;
          addr[63] = loop_63[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_64 = 1'b0;
        addr[64] = 3'b0;
        for (loop_64 = 0; loop_64 < NUM_CELL; loop_64++) begin
         if ({b[0],a[2]}) == loop_64[1:0]) begin
          match_flag_64 = 1'b1;
          addr[64] = loop_64[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_65 = 1'b0;
        addr[65] = 3'b0;
        for (loop_65 = 0; loop_65 < NUM_CELL; loop_65++) begin
         if ({b[1],a[2]}) == loop_65[1:0]) begin
          match_flag_65 = 1'b1;
          addr[65] = loop_65[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_66 = 1'b0;
        addr[66] = 3'b0;
        for (loop_66 = 0; loop_66 < NUM_CELL; loop_66++) begin
         if ({b[2],a[2]}) == loop_66[1:0]) begin
          match_flag_66 = 1'b1;
          addr[66] = loop_66[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_67 = 1'b0;
        addr[67] = 3'b0;
        for (loop_67 = 0; loop_67 < NUM_CELL; loop_67++) begin
         if ({b[3],a[2]}) == loop_67[1:0]) begin
          match_flag_67 = 1'b1;
          addr[67] = loop_67[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_68 = 1'b0;
        addr[68] = 3'b0;
        for (loop_68 = 0; loop_68 < NUM_CELL; loop_68++) begin
         if ({b[4],a[2]}) == loop_68[1:0]) begin
          match_flag_68 = 1'b1;
          addr[68] = loop_68[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_69 = 1'b0;
        addr[69] = 3'b0;
        for (loop_69 = 0; loop_69 < NUM_CELL; loop_69++) begin
         if ({b[5],a[2]}) == loop_69[1:0]) begin
          match_flag_69 = 1'b1;
          addr[69] = loop_69[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_70 = 1'b0;
        addr[70] = 3'b0;
        for (loop_70 = 0; loop_70 < NUM_CELL; loop_70++) begin
         if ({b[6],a[2]}) == loop_70[1:0]) begin
          match_flag_70 = 1'b1;
          addr[70] = loop_70[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_71 = 1'b0;
        addr[71] = 3'b0;
        for (loop_71 = 0; loop_71 < NUM_CELL; loop_71++) begin
         if ({b[7],a[2]}) == loop_71[1:0]) begin
          match_flag_71 = 1'b1;
          addr[71] = loop_71[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_72 = 1'b0;
        addr[72] = 3'b0;
        for (loop_72 = 0; loop_72 < NUM_CELL; loop_72++) begin
         if ({b[8],a[2]}) == loop_72[1:0]) begin
          match_flag_72 = 1'b1;
          addr[72] = loop_72[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_73 = 1'b0;
        addr[73] = 3'b0;
        for (loop_73 = 0; loop_73 < NUM_CELL; loop_73++) begin
         if ({b[9],a[2]}) == loop_73[1:0]) begin
          match_flag_73 = 1'b1;
          addr[73] = loop_73[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_74 = 1'b0;
        addr[74] = 3'b0;
        for (loop_74 = 0; loop_74 < NUM_CELL; loop_74++) begin
         if ({b[10],a[2]}) == loop_74[1:0]) begin
          match_flag_74 = 1'b1;
          addr[74] = loop_74[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_75 = 1'b0;
        addr[75] = 3'b0;
        for (loop_75 = 0; loop_75 < NUM_CELL; loop_75++) begin
         if ({b[11],a[2]}) == loop_75[1:0]) begin
          match_flag_75 = 1'b1;
          addr[75] = loop_75[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_76 = 1'b0;
        addr[76] = 3'b0;
        for (loop_76 = 0; loop_76 < NUM_CELL; loop_76++) begin
         if ({b[12],a[2]}) == loop_76[1:0]) begin
          match_flag_76 = 1'b1;
          addr[76] = loop_76[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_77 = 1'b0;
        addr[77] = 3'b0;
        for (loop_77 = 0; loop_77 < NUM_CELL; loop_77++) begin
         if ({b[13],a[2]}) == loop_77[1:0]) begin
          match_flag_77 = 1'b1;
          addr[77] = loop_77[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_78 = 1'b0;
        addr[78] = 3'b0;
        for (loop_78 = 0; loop_78 < NUM_CELL; loop_78++) begin
         if ({b[14],a[2]}) == loop_78[1:0]) begin
          match_flag_78 = 1'b1;
          addr[78] = loop_78[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_79 = 1'b0;
        addr[79] = 3'b0;
        for (loop_79 = 0; loop_79 < NUM_CELL; loop_79++) begin
         if ({b[15],a[2]}) == loop_79[1:0]) begin
          match_flag_79 = 1'b1;
          addr[79] = loop_79[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_80 = 1'b0;
        addr[80] = 3'b0;
        for (loop_80 = 0; loop_80 < NUM_CELL; loop_80++) begin
         if ({b[16],a[2]}) == loop_80[1:0]) begin
          match_flag_80 = 1'b1;
          addr[80] = loop_80[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_81 = 1'b0;
        addr[81] = 3'b0;
        for (loop_81 = 0; loop_81 < NUM_CELL; loop_81++) begin
         if ({b[17],a[2]}) == loop_81[1:0]) begin
          match_flag_81 = 1'b1;
          addr[81] = loop_81[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_82 = 1'b0;
        addr[82] = 3'b0;
        for (loop_82 = 0; loop_82 < NUM_CELL; loop_82++) begin
         if ({b[18],a[2]}) == loop_82[1:0]) begin
          match_flag_82 = 1'b1;
          addr[82] = loop_82[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_83 = 1'b0;
        addr[83] = 3'b0;
        for (loop_83 = 0; loop_83 < NUM_CELL; loop_83++) begin
         if ({b[19],a[2]}) == loop_83[1:0]) begin
          match_flag_83 = 1'b1;
          addr[83] = loop_83[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_84 = 1'b0;
        addr[84] = 3'b0;
        for (loop_84 = 0; loop_84 < NUM_CELL; loop_84++) begin
         if ({b[20],a[2]}) == loop_84[1:0]) begin
          match_flag_84 = 1'b1;
          addr[84] = loop_84[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_85 = 1'b0;
        addr[85] = 3'b0;
        for (loop_85 = 0; loop_85 < NUM_CELL; loop_85++) begin
         if ({b[21],a[2]}) == loop_85[1:0]) begin
          match_flag_85 = 1'b1;
          addr[85] = loop_85[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_86 = 1'b0;
        addr[86] = 3'b0;
        for (loop_86 = 0; loop_86 < NUM_CELL; loop_86++) begin
         if ({b[22],a[2]}) == loop_86[1:0]) begin
          match_flag_86 = 1'b1;
          addr[86] = loop_86[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_87 = 1'b0;
        addr[87] = 3'b0;
        for (loop_87 = 0; loop_87 < NUM_CELL; loop_87++) begin
         if ({b[23],a[2]}) == loop_87[1:0]) begin
          match_flag_87 = 1'b1;
          addr[87] = loop_87[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_88 = 1'b0;
        addr[88] = 3'b0;
        for (loop_88 = 0; loop_88 < NUM_CELL; loop_88++) begin
         if ({b[24],a[2]}) == loop_88[1:0]) begin
          match_flag_88 = 1'b1;
          addr[88] = loop_88[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_89 = 1'b0;
        addr[89] = 3'b0;
        for (loop_89 = 0; loop_89 < NUM_CELL; loop_89++) begin
         if ({b[25],a[2]}) == loop_89[1:0]) begin
          match_flag_89 = 1'b1;
          addr[89] = loop_89[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_90 = 1'b0;
        addr[90] = 3'b0;
        for (loop_90 = 0; loop_90 < NUM_CELL; loop_90++) begin
         if ({b[26],a[2]}) == loop_90[1:0]) begin
          match_flag_90 = 1'b1;
          addr[90] = loop_90[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_91 = 1'b0;
        addr[91] = 3'b0;
        for (loop_91 = 0; loop_91 < NUM_CELL; loop_91++) begin
         if ({b[27],a[2]}) == loop_91[1:0]) begin
          match_flag_91 = 1'b1;
          addr[91] = loop_91[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_92 = 1'b0;
        addr[92] = 3'b0;
        for (loop_92 = 0; loop_92 < NUM_CELL; loop_92++) begin
         if ({b[28],a[2]}) == loop_92[1:0]) begin
          match_flag_92 = 1'b1;
          addr[92] = loop_92[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_93 = 1'b0;
        addr[93] = 3'b0;
        for (loop_93 = 0; loop_93 < NUM_CELL; loop_93++) begin
         if ({b[29],a[2]}) == loop_93[1:0]) begin
          match_flag_93 = 1'b1;
          addr[93] = loop_93[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_94 = 1'b0;
        addr[94] = 3'b0;
        for (loop_94 = 0; loop_94 < NUM_CELL; loop_94++) begin
         if ({b[30],a[2]}) == loop_94[1:0]) begin
          match_flag_94 = 1'b1;
          addr[94] = loop_94[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_95 = 1'b0;
        addr[95] = 3'b0;
        for (loop_95 = 0; loop_95 < NUM_CELL; loop_95++) begin
         if ({b[31],a[2]}) == loop_95[1:0]) begin
          match_flag_95 = 1'b1;
          addr[95] = loop_95[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_96 = 1'b0;
        addr[96] = 3'b0;
        for (loop_96 = 0; loop_96 < NUM_CELL; loop_96++) begin
         if ({b[0],a[3]}) == loop_96[1:0]) begin
          match_flag_96 = 1'b1;
          addr[96] = loop_96[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_97 = 1'b0;
        addr[97] = 3'b0;
        for (loop_97 = 0; loop_97 < NUM_CELL; loop_97++) begin
         if ({b[1],a[3]}) == loop_97[1:0]) begin
          match_flag_97 = 1'b1;
          addr[97] = loop_97[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_98 = 1'b0;
        addr[98] = 3'b0;
        for (loop_98 = 0; loop_98 < NUM_CELL; loop_98++) begin
         if ({b[2],a[3]}) == loop_98[1:0]) begin
          match_flag_98 = 1'b1;
          addr[98] = loop_98[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_99 = 1'b0;
        addr[99] = 3'b0;
        for (loop_99 = 0; loop_99 < NUM_CELL; loop_99++) begin
         if ({b[3],a[3]}) == loop_99[1:0]) begin
          match_flag_99 = 1'b1;
          addr[99] = loop_99[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_100 = 1'b0;
        addr[100] = 3'b0;
        for (loop_100 = 0; loop_100 < NUM_CELL; loop_100++) begin
         if ({b[4],a[3]}) == loop_100[1:0]) begin
          match_flag_100 = 1'b1;
          addr[100] = loop_100[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_101 = 1'b0;
        addr[101] = 3'b0;
        for (loop_101 = 0; loop_101 < NUM_CELL; loop_101++) begin
         if ({b[5],a[3]}) == loop_101[1:0]) begin
          match_flag_101 = 1'b1;
          addr[101] = loop_101[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_102 = 1'b0;
        addr[102] = 3'b0;
        for (loop_102 = 0; loop_102 < NUM_CELL; loop_102++) begin
         if ({b[6],a[3]}) == loop_102[1:0]) begin
          match_flag_102 = 1'b1;
          addr[102] = loop_102[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_103 = 1'b0;
        addr[103] = 3'b0;
        for (loop_103 = 0; loop_103 < NUM_CELL; loop_103++) begin
         if ({b[7],a[3]}) == loop_103[1:0]) begin
          match_flag_103 = 1'b1;
          addr[103] = loop_103[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_104 = 1'b0;
        addr[104] = 3'b0;
        for (loop_104 = 0; loop_104 < NUM_CELL; loop_104++) begin
         if ({b[8],a[3]}) == loop_104[1:0]) begin
          match_flag_104 = 1'b1;
          addr[104] = loop_104[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_105 = 1'b0;
        addr[105] = 3'b0;
        for (loop_105 = 0; loop_105 < NUM_CELL; loop_105++) begin
         if ({b[9],a[3]}) == loop_105[1:0]) begin
          match_flag_105 = 1'b1;
          addr[105] = loop_105[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_106 = 1'b0;
        addr[106] = 3'b0;
        for (loop_106 = 0; loop_106 < NUM_CELL; loop_106++) begin
         if ({b[10],a[3]}) == loop_106[1:0]) begin
          match_flag_106 = 1'b1;
          addr[106] = loop_106[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_107 = 1'b0;
        addr[107] = 3'b0;
        for (loop_107 = 0; loop_107 < NUM_CELL; loop_107++) begin
         if ({b[11],a[3]}) == loop_107[1:0]) begin
          match_flag_107 = 1'b1;
          addr[107] = loop_107[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_108 = 1'b0;
        addr[108] = 3'b0;
        for (loop_108 = 0; loop_108 < NUM_CELL; loop_108++) begin
         if ({b[12],a[3]}) == loop_108[1:0]) begin
          match_flag_108 = 1'b1;
          addr[108] = loop_108[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_109 = 1'b0;
        addr[109] = 3'b0;
        for (loop_109 = 0; loop_109 < NUM_CELL; loop_109++) begin
         if ({b[13],a[3]}) == loop_109[1:0]) begin
          match_flag_109 = 1'b1;
          addr[109] = loop_109[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_110 = 1'b0;
        addr[110] = 3'b0;
        for (loop_110 = 0; loop_110 < NUM_CELL; loop_110++) begin
         if ({b[14],a[3]}) == loop_110[1:0]) begin
          match_flag_110 = 1'b1;
          addr[110] = loop_110[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_111 = 1'b0;
        addr[111] = 3'b0;
        for (loop_111 = 0; loop_111 < NUM_CELL; loop_111++) begin
         if ({b[15],a[3]}) == loop_111[1:0]) begin
          match_flag_111 = 1'b1;
          addr[111] = loop_111[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_112 = 1'b0;
        addr[112] = 3'b0;
        for (loop_112 = 0; loop_112 < NUM_CELL; loop_112++) begin
         if ({b[16],a[3]}) == loop_112[1:0]) begin
          match_flag_112 = 1'b1;
          addr[112] = loop_112[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_113 = 1'b0;
        addr[113] = 3'b0;
        for (loop_113 = 0; loop_113 < NUM_CELL; loop_113++) begin
         if ({b[17],a[3]}) == loop_113[1:0]) begin
          match_flag_113 = 1'b1;
          addr[113] = loop_113[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_114 = 1'b0;
        addr[114] = 3'b0;
        for (loop_114 = 0; loop_114 < NUM_CELL; loop_114++) begin
         if ({b[18],a[3]}) == loop_114[1:0]) begin
          match_flag_114 = 1'b1;
          addr[114] = loop_114[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_115 = 1'b0;
        addr[115] = 3'b0;
        for (loop_115 = 0; loop_115 < NUM_CELL; loop_115++) begin
         if ({b[19],a[3]}) == loop_115[1:0]) begin
          match_flag_115 = 1'b1;
          addr[115] = loop_115[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_116 = 1'b0;
        addr[116] = 3'b0;
        for (loop_116 = 0; loop_116 < NUM_CELL; loop_116++) begin
         if ({b[20],a[3]}) == loop_116[1:0]) begin
          match_flag_116 = 1'b1;
          addr[116] = loop_116[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_117 = 1'b0;
        addr[117] = 3'b0;
        for (loop_117 = 0; loop_117 < NUM_CELL; loop_117++) begin
         if ({b[21],a[3]}) == loop_117[1:0]) begin
          match_flag_117 = 1'b1;
          addr[117] = loop_117[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_118 = 1'b0;
        addr[118] = 3'b0;
        for (loop_118 = 0; loop_118 < NUM_CELL; loop_118++) begin
         if ({b[22],a[3]}) == loop_118[1:0]) begin
          match_flag_118 = 1'b1;
          addr[118] = loop_118[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_119 = 1'b0;
        addr[119] = 3'b0;
        for (loop_119 = 0; loop_119 < NUM_CELL; loop_119++) begin
         if ({b[23],a[3]}) == loop_119[1:0]) begin
          match_flag_119 = 1'b1;
          addr[119] = loop_119[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_120 = 1'b0;
        addr[120] = 3'b0;
        for (loop_120 = 0; loop_120 < NUM_CELL; loop_120++) begin
         if ({b[24],a[3]}) == loop_120[1:0]) begin
          match_flag_120 = 1'b1;
          addr[120] = loop_120[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_121 = 1'b0;
        addr[121] = 3'b0;
        for (loop_121 = 0; loop_121 < NUM_CELL; loop_121++) begin
         if ({b[25],a[3]}) == loop_121[1:0]) begin
          match_flag_121 = 1'b1;
          addr[121] = loop_121[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_122 = 1'b0;
        addr[122] = 3'b0;
        for (loop_122 = 0; loop_122 < NUM_CELL; loop_122++) begin
         if ({b[26],a[3]}) == loop_122[1:0]) begin
          match_flag_122 = 1'b1;
          addr[122] = loop_122[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_123 = 1'b0;
        addr[123] = 3'b0;
        for (loop_123 = 0; loop_123 < NUM_CELL; loop_123++) begin
         if ({b[27],a[3]}) == loop_123[1:0]) begin
          match_flag_123 = 1'b1;
          addr[123] = loop_123[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_124 = 1'b0;
        addr[124] = 3'b0;
        for (loop_124 = 0; loop_124 < NUM_CELL; loop_124++) begin
         if ({b[28],a[3]}) == loop_124[1:0]) begin
          match_flag_124 = 1'b1;
          addr[124] = loop_124[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_125 = 1'b0;
        addr[125] = 3'b0;
        for (loop_125 = 0; loop_125 < NUM_CELL; loop_125++) begin
         if ({b[29],a[3]}) == loop_125[1:0]) begin
          match_flag_125 = 1'b1;
          addr[125] = loop_125[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_126 = 1'b0;
        addr[126] = 3'b0;
        for (loop_126 = 0; loop_126 < NUM_CELL; loop_126++) begin
         if ({b[30],a[3]}) == loop_126[1:0]) begin
          match_flag_126 = 1'b1;
          addr[126] = loop_126[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_127 = 1'b0;
        addr[127] = 3'b0;
        for (loop_127 = 0; loop_127 < NUM_CELL; loop_127++) begin
         if ({b[31],a[3]}) == loop_127[1:0]) begin
          match_flag_127 = 1'b1;
          addr[127] = loop_127[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_128 = 1'b0;
        addr[128] = 3'b0;
        for (loop_128 = 0; loop_128 < NUM_CELL; loop_128++) begin
         if ({b[0],a[4]}) == loop_128[1:0]) begin
          match_flag_128 = 1'b1;
          addr[128] = loop_128[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_129 = 1'b0;
        addr[129] = 3'b0;
        for (loop_129 = 0; loop_129 < NUM_CELL; loop_129++) begin
         if ({b[1],a[4]}) == loop_129[1:0]) begin
          match_flag_129 = 1'b1;
          addr[129] = loop_129[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_130 = 1'b0;
        addr[130] = 3'b0;
        for (loop_130 = 0; loop_130 < NUM_CELL; loop_130++) begin
         if ({b[2],a[4]}) == loop_130[1:0]) begin
          match_flag_130 = 1'b1;
          addr[130] = loop_130[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_131 = 1'b0;
        addr[131] = 3'b0;
        for (loop_131 = 0; loop_131 < NUM_CELL; loop_131++) begin
         if ({b[3],a[4]}) == loop_131[1:0]) begin
          match_flag_131 = 1'b1;
          addr[131] = loop_131[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_132 = 1'b0;
        addr[132] = 3'b0;
        for (loop_132 = 0; loop_132 < NUM_CELL; loop_132++) begin
         if ({b[4],a[4]}) == loop_132[1:0]) begin
          match_flag_132 = 1'b1;
          addr[132] = loop_132[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_133 = 1'b0;
        addr[133] = 3'b0;
        for (loop_133 = 0; loop_133 < NUM_CELL; loop_133++) begin
         if ({b[5],a[4]}) == loop_133[1:0]) begin
          match_flag_133 = 1'b1;
          addr[133] = loop_133[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_134 = 1'b0;
        addr[134] = 3'b0;
        for (loop_134 = 0; loop_134 < NUM_CELL; loop_134++) begin
         if ({b[6],a[4]}) == loop_134[1:0]) begin
          match_flag_134 = 1'b1;
          addr[134] = loop_134[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_135 = 1'b0;
        addr[135] = 3'b0;
        for (loop_135 = 0; loop_135 < NUM_CELL; loop_135++) begin
         if ({b[7],a[4]}) == loop_135[1:0]) begin
          match_flag_135 = 1'b1;
          addr[135] = loop_135[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_136 = 1'b0;
        addr[136] = 3'b0;
        for (loop_136 = 0; loop_136 < NUM_CELL; loop_136++) begin
         if ({b[8],a[4]}) == loop_136[1:0]) begin
          match_flag_136 = 1'b1;
          addr[136] = loop_136[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_137 = 1'b0;
        addr[137] = 3'b0;
        for (loop_137 = 0; loop_137 < NUM_CELL; loop_137++) begin
         if ({b[9],a[4]}) == loop_137[1:0]) begin
          match_flag_137 = 1'b1;
          addr[137] = loop_137[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_138 = 1'b0;
        addr[138] = 3'b0;
        for (loop_138 = 0; loop_138 < NUM_CELL; loop_138++) begin
         if ({b[10],a[4]}) == loop_138[1:0]) begin
          match_flag_138 = 1'b1;
          addr[138] = loop_138[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_139 = 1'b0;
        addr[139] = 3'b0;
        for (loop_139 = 0; loop_139 < NUM_CELL; loop_139++) begin
         if ({b[11],a[4]}) == loop_139[1:0]) begin
          match_flag_139 = 1'b1;
          addr[139] = loop_139[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_140 = 1'b0;
        addr[140] = 3'b0;
        for (loop_140 = 0; loop_140 < NUM_CELL; loop_140++) begin
         if ({b[12],a[4]}) == loop_140[1:0]) begin
          match_flag_140 = 1'b1;
          addr[140] = loop_140[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_141 = 1'b0;
        addr[141] = 3'b0;
        for (loop_141 = 0; loop_141 < NUM_CELL; loop_141++) begin
         if ({b[13],a[4]}) == loop_141[1:0]) begin
          match_flag_141 = 1'b1;
          addr[141] = loop_141[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_142 = 1'b0;
        addr[142] = 3'b0;
        for (loop_142 = 0; loop_142 < NUM_CELL; loop_142++) begin
         if ({b[14],a[4]}) == loop_142[1:0]) begin
          match_flag_142 = 1'b1;
          addr[142] = loop_142[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_143 = 1'b0;
        addr[143] = 3'b0;
        for (loop_143 = 0; loop_143 < NUM_CELL; loop_143++) begin
         if ({b[15],a[4]}) == loop_143[1:0]) begin
          match_flag_143 = 1'b1;
          addr[143] = loop_143[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_144 = 1'b0;
        addr[144] = 3'b0;
        for (loop_144 = 0; loop_144 < NUM_CELL; loop_144++) begin
         if ({b[16],a[4]}) == loop_144[1:0]) begin
          match_flag_144 = 1'b1;
          addr[144] = loop_144[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_145 = 1'b0;
        addr[145] = 3'b0;
        for (loop_145 = 0; loop_145 < NUM_CELL; loop_145++) begin
         if ({b[17],a[4]}) == loop_145[1:0]) begin
          match_flag_145 = 1'b1;
          addr[145] = loop_145[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_146 = 1'b0;
        addr[146] = 3'b0;
        for (loop_146 = 0; loop_146 < NUM_CELL; loop_146++) begin
         if ({b[18],a[4]}) == loop_146[1:0]) begin
          match_flag_146 = 1'b1;
          addr[146] = loop_146[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_147 = 1'b0;
        addr[147] = 3'b0;
        for (loop_147 = 0; loop_147 < NUM_CELL; loop_147++) begin
         if ({b[19],a[4]}) == loop_147[1:0]) begin
          match_flag_147 = 1'b1;
          addr[147] = loop_147[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_148 = 1'b0;
        addr[148] = 3'b0;
        for (loop_148 = 0; loop_148 < NUM_CELL; loop_148++) begin
         if ({b[20],a[4]}) == loop_148[1:0]) begin
          match_flag_148 = 1'b1;
          addr[148] = loop_148[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_149 = 1'b0;
        addr[149] = 3'b0;
        for (loop_149 = 0; loop_149 < NUM_CELL; loop_149++) begin
         if ({b[21],a[4]}) == loop_149[1:0]) begin
          match_flag_149 = 1'b1;
          addr[149] = loop_149[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_150 = 1'b0;
        addr[150] = 3'b0;
        for (loop_150 = 0; loop_150 < NUM_CELL; loop_150++) begin
         if ({b[22],a[4]}) == loop_150[1:0]) begin
          match_flag_150 = 1'b1;
          addr[150] = loop_150[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_151 = 1'b0;
        addr[151] = 3'b0;
        for (loop_151 = 0; loop_151 < NUM_CELL; loop_151++) begin
         if ({b[23],a[4]}) == loop_151[1:0]) begin
          match_flag_151 = 1'b1;
          addr[151] = loop_151[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_152 = 1'b0;
        addr[152] = 3'b0;
        for (loop_152 = 0; loop_152 < NUM_CELL; loop_152++) begin
         if ({b[24],a[4]}) == loop_152[1:0]) begin
          match_flag_152 = 1'b1;
          addr[152] = loop_152[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_153 = 1'b0;
        addr[153] = 3'b0;
        for (loop_153 = 0; loop_153 < NUM_CELL; loop_153++) begin
         if ({b[25],a[4]}) == loop_153[1:0]) begin
          match_flag_153 = 1'b1;
          addr[153] = loop_153[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_154 = 1'b0;
        addr[154] = 3'b0;
        for (loop_154 = 0; loop_154 < NUM_CELL; loop_154++) begin
         if ({b[26],a[4]}) == loop_154[1:0]) begin
          match_flag_154 = 1'b1;
          addr[154] = loop_154[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_155 = 1'b0;
        addr[155] = 3'b0;
        for (loop_155 = 0; loop_155 < NUM_CELL; loop_155++) begin
         if ({b[27],a[4]}) == loop_155[1:0]) begin
          match_flag_155 = 1'b1;
          addr[155] = loop_155[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_156 = 1'b0;
        addr[156] = 3'b0;
        for (loop_156 = 0; loop_156 < NUM_CELL; loop_156++) begin
         if ({b[28],a[4]}) == loop_156[1:0]) begin
          match_flag_156 = 1'b1;
          addr[156] = loop_156[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_157 = 1'b0;
        addr[157] = 3'b0;
        for (loop_157 = 0; loop_157 < NUM_CELL; loop_157++) begin
         if ({b[29],a[4]}) == loop_157[1:0]) begin
          match_flag_157 = 1'b1;
          addr[157] = loop_157[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_158 = 1'b0;
        addr[158] = 3'b0;
        for (loop_158 = 0; loop_158 < NUM_CELL; loop_158++) begin
         if ({b[30],a[4]}) == loop_158[1:0]) begin
          match_flag_158 = 1'b1;
          addr[158] = loop_158[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_159 = 1'b0;
        addr[159] = 3'b0;
        for (loop_159 = 0; loop_159 < NUM_CELL; loop_159++) begin
         if ({b[31],a[4]}) == loop_159[1:0]) begin
          match_flag_159 = 1'b1;
          addr[159] = loop_159[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_160 = 1'b0;
        addr[160] = 3'b0;
        for (loop_160 = 0; loop_160 < NUM_CELL; loop_160++) begin
         if ({b[0],a[5]}) == loop_160[1:0]) begin
          match_flag_160 = 1'b1;
          addr[160] = loop_160[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_161 = 1'b0;
        addr[161] = 3'b0;
        for (loop_161 = 0; loop_161 < NUM_CELL; loop_161++) begin
         if ({b[1],a[5]}) == loop_161[1:0]) begin
          match_flag_161 = 1'b1;
          addr[161] = loop_161[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_162 = 1'b0;
        addr[162] = 3'b0;
        for (loop_162 = 0; loop_162 < NUM_CELL; loop_162++) begin
         if ({b[2],a[5]}) == loop_162[1:0]) begin
          match_flag_162 = 1'b1;
          addr[162] = loop_162[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_163 = 1'b0;
        addr[163] = 3'b0;
        for (loop_163 = 0; loop_163 < NUM_CELL; loop_163++) begin
         if ({b[3],a[5]}) == loop_163[1:0]) begin
          match_flag_163 = 1'b1;
          addr[163] = loop_163[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_164 = 1'b0;
        addr[164] = 3'b0;
        for (loop_164 = 0; loop_164 < NUM_CELL; loop_164++) begin
         if ({b[4],a[5]}) == loop_164[1:0]) begin
          match_flag_164 = 1'b1;
          addr[164] = loop_164[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_165 = 1'b0;
        addr[165] = 3'b0;
        for (loop_165 = 0; loop_165 < NUM_CELL; loop_165++) begin
         if ({b[5],a[5]}) == loop_165[1:0]) begin
          match_flag_165 = 1'b1;
          addr[165] = loop_165[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_166 = 1'b0;
        addr[166] = 3'b0;
        for (loop_166 = 0; loop_166 < NUM_CELL; loop_166++) begin
         if ({b[6],a[5]}) == loop_166[1:0]) begin
          match_flag_166 = 1'b1;
          addr[166] = loop_166[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_167 = 1'b0;
        addr[167] = 3'b0;
        for (loop_167 = 0; loop_167 < NUM_CELL; loop_167++) begin
         if ({b[7],a[5]}) == loop_167[1:0]) begin
          match_flag_167 = 1'b1;
          addr[167] = loop_167[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_168 = 1'b0;
        addr[168] = 3'b0;
        for (loop_168 = 0; loop_168 < NUM_CELL; loop_168++) begin
         if ({b[8],a[5]}) == loop_168[1:0]) begin
          match_flag_168 = 1'b1;
          addr[168] = loop_168[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_169 = 1'b0;
        addr[169] = 3'b0;
        for (loop_169 = 0; loop_169 < NUM_CELL; loop_169++) begin
         if ({b[9],a[5]}) == loop_169[1:0]) begin
          match_flag_169 = 1'b1;
          addr[169] = loop_169[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_170 = 1'b0;
        addr[170] = 3'b0;
        for (loop_170 = 0; loop_170 < NUM_CELL; loop_170++) begin
         if ({b[10],a[5]}) == loop_170[1:0]) begin
          match_flag_170 = 1'b1;
          addr[170] = loop_170[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_171 = 1'b0;
        addr[171] = 3'b0;
        for (loop_171 = 0; loop_171 < NUM_CELL; loop_171++) begin
         if ({b[11],a[5]}) == loop_171[1:0]) begin
          match_flag_171 = 1'b1;
          addr[171] = loop_171[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_172 = 1'b0;
        addr[172] = 3'b0;
        for (loop_172 = 0; loop_172 < NUM_CELL; loop_172++) begin
         if ({b[12],a[5]}) == loop_172[1:0]) begin
          match_flag_172 = 1'b1;
          addr[172] = loop_172[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_173 = 1'b0;
        addr[173] = 3'b0;
        for (loop_173 = 0; loop_173 < NUM_CELL; loop_173++) begin
         if ({b[13],a[5]}) == loop_173[1:0]) begin
          match_flag_173 = 1'b1;
          addr[173] = loop_173[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_174 = 1'b0;
        addr[174] = 3'b0;
        for (loop_174 = 0; loop_174 < NUM_CELL; loop_174++) begin
         if ({b[14],a[5]}) == loop_174[1:0]) begin
          match_flag_174 = 1'b1;
          addr[174] = loop_174[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_175 = 1'b0;
        addr[175] = 3'b0;
        for (loop_175 = 0; loop_175 < NUM_CELL; loop_175++) begin
         if ({b[15],a[5]}) == loop_175[1:0]) begin
          match_flag_175 = 1'b1;
          addr[175] = loop_175[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_176 = 1'b0;
        addr[176] = 3'b0;
        for (loop_176 = 0; loop_176 < NUM_CELL; loop_176++) begin
         if ({b[16],a[5]}) == loop_176[1:0]) begin
          match_flag_176 = 1'b1;
          addr[176] = loop_176[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_177 = 1'b0;
        addr[177] = 3'b0;
        for (loop_177 = 0; loop_177 < NUM_CELL; loop_177++) begin
         if ({b[17],a[5]}) == loop_177[1:0]) begin
          match_flag_177 = 1'b1;
          addr[177] = loop_177[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_178 = 1'b0;
        addr[178] = 3'b0;
        for (loop_178 = 0; loop_178 < NUM_CELL; loop_178++) begin
         if ({b[18],a[5]}) == loop_178[1:0]) begin
          match_flag_178 = 1'b1;
          addr[178] = loop_178[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_179 = 1'b0;
        addr[179] = 3'b0;
        for (loop_179 = 0; loop_179 < NUM_CELL; loop_179++) begin
         if ({b[19],a[5]}) == loop_179[1:0]) begin
          match_flag_179 = 1'b1;
          addr[179] = loop_179[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_180 = 1'b0;
        addr[180] = 3'b0;
        for (loop_180 = 0; loop_180 < NUM_CELL; loop_180++) begin
         if ({b[20],a[5]}) == loop_180[1:0]) begin
          match_flag_180 = 1'b1;
          addr[180] = loop_180[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_181 = 1'b0;
        addr[181] = 3'b0;
        for (loop_181 = 0; loop_181 < NUM_CELL; loop_181++) begin
         if ({b[21],a[5]}) == loop_181[1:0]) begin
          match_flag_181 = 1'b1;
          addr[181] = loop_181[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_182 = 1'b0;
        addr[182] = 3'b0;
        for (loop_182 = 0; loop_182 < NUM_CELL; loop_182++) begin
         if ({b[22],a[5]}) == loop_182[1:0]) begin
          match_flag_182 = 1'b1;
          addr[182] = loop_182[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_183 = 1'b0;
        addr[183] = 3'b0;
        for (loop_183 = 0; loop_183 < NUM_CELL; loop_183++) begin
         if ({b[23],a[5]}) == loop_183[1:0]) begin
          match_flag_183 = 1'b1;
          addr[183] = loop_183[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_184 = 1'b0;
        addr[184] = 3'b0;
        for (loop_184 = 0; loop_184 < NUM_CELL; loop_184++) begin
         if ({b[24],a[5]}) == loop_184[1:0]) begin
          match_flag_184 = 1'b1;
          addr[184] = loop_184[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_185 = 1'b0;
        addr[185] = 3'b0;
        for (loop_185 = 0; loop_185 < NUM_CELL; loop_185++) begin
         if ({b[25],a[5]}) == loop_185[1:0]) begin
          match_flag_185 = 1'b1;
          addr[185] = loop_185[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_186 = 1'b0;
        addr[186] = 3'b0;
        for (loop_186 = 0; loop_186 < NUM_CELL; loop_186++) begin
         if ({b[26],a[5]}) == loop_186[1:0]) begin
          match_flag_186 = 1'b1;
          addr[186] = loop_186[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_187 = 1'b0;
        addr[187] = 3'b0;
        for (loop_187 = 0; loop_187 < NUM_CELL; loop_187++) begin
         if ({b[27],a[5]}) == loop_187[1:0]) begin
          match_flag_187 = 1'b1;
          addr[187] = loop_187[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_188 = 1'b0;
        addr[188] = 3'b0;
        for (loop_188 = 0; loop_188 < NUM_CELL; loop_188++) begin
         if ({b[28],a[5]}) == loop_188[1:0]) begin
          match_flag_188 = 1'b1;
          addr[188] = loop_188[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_189 = 1'b0;
        addr[189] = 3'b0;
        for (loop_189 = 0; loop_189 < NUM_CELL; loop_189++) begin
         if ({b[29],a[5]}) == loop_189[1:0]) begin
          match_flag_189 = 1'b1;
          addr[189] = loop_189[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_190 = 1'b0;
        addr[190] = 3'b0;
        for (loop_190 = 0; loop_190 < NUM_CELL; loop_190++) begin
         if ({b[30],a[5]}) == loop_190[1:0]) begin
          match_flag_190 = 1'b1;
          addr[190] = loop_190[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_191 = 1'b0;
        addr[191] = 3'b0;
        for (loop_191 = 0; loop_191 < NUM_CELL; loop_191++) begin
         if ({b[31],a[5]}) == loop_191[1:0]) begin
          match_flag_191 = 1'b1;
          addr[191] = loop_191[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_192 = 1'b0;
        addr[192] = 3'b0;
        for (loop_192 = 0; loop_192 < NUM_CELL; loop_192++) begin
         if ({b[0],a[6]}) == loop_192[1:0]) begin
          match_flag_192 = 1'b1;
          addr[192] = loop_192[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_193 = 1'b0;
        addr[193] = 3'b0;
        for (loop_193 = 0; loop_193 < NUM_CELL; loop_193++) begin
         if ({b[1],a[6]}) == loop_193[1:0]) begin
          match_flag_193 = 1'b1;
          addr[193] = loop_193[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_194 = 1'b0;
        addr[194] = 3'b0;
        for (loop_194 = 0; loop_194 < NUM_CELL; loop_194++) begin
         if ({b[2],a[6]}) == loop_194[1:0]) begin
          match_flag_194 = 1'b1;
          addr[194] = loop_194[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_195 = 1'b0;
        addr[195] = 3'b0;
        for (loop_195 = 0; loop_195 < NUM_CELL; loop_195++) begin
         if ({b[3],a[6]}) == loop_195[1:0]) begin
          match_flag_195 = 1'b1;
          addr[195] = loop_195[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_196 = 1'b0;
        addr[196] = 3'b0;
        for (loop_196 = 0; loop_196 < NUM_CELL; loop_196++) begin
         if ({b[4],a[6]}) == loop_196[1:0]) begin
          match_flag_196 = 1'b1;
          addr[196] = loop_196[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_197 = 1'b0;
        addr[197] = 3'b0;
        for (loop_197 = 0; loop_197 < NUM_CELL; loop_197++) begin
         if ({b[5],a[6]}) == loop_197[1:0]) begin
          match_flag_197 = 1'b1;
          addr[197] = loop_197[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_198 = 1'b0;
        addr[198] = 3'b0;
        for (loop_198 = 0; loop_198 < NUM_CELL; loop_198++) begin
         if ({b[6],a[6]}) == loop_198[1:0]) begin
          match_flag_198 = 1'b1;
          addr[198] = loop_198[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_199 = 1'b0;
        addr[199] = 3'b0;
        for (loop_199 = 0; loop_199 < NUM_CELL; loop_199++) begin
         if ({b[7],a[6]}) == loop_199[1:0]) begin
          match_flag_199 = 1'b1;
          addr[199] = loop_199[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_200 = 1'b0;
        addr[200] = 3'b0;
        for (loop_200 = 0; loop_200 < NUM_CELL; loop_200++) begin
         if ({b[8],a[6]}) == loop_200[1:0]) begin
          match_flag_200 = 1'b1;
          addr[200] = loop_200[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_201 = 1'b0;
        addr[201] = 3'b0;
        for (loop_201 = 0; loop_201 < NUM_CELL; loop_201++) begin
         if ({b[9],a[6]}) == loop_201[1:0]) begin
          match_flag_201 = 1'b1;
          addr[201] = loop_201[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_202 = 1'b0;
        addr[202] = 3'b0;
        for (loop_202 = 0; loop_202 < NUM_CELL; loop_202++) begin
         if ({b[10],a[6]}) == loop_202[1:0]) begin
          match_flag_202 = 1'b1;
          addr[202] = loop_202[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_203 = 1'b0;
        addr[203] = 3'b0;
        for (loop_203 = 0; loop_203 < NUM_CELL; loop_203++) begin
         if ({b[11],a[6]}) == loop_203[1:0]) begin
          match_flag_203 = 1'b1;
          addr[203] = loop_203[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_204 = 1'b0;
        addr[204] = 3'b0;
        for (loop_204 = 0; loop_204 < NUM_CELL; loop_204++) begin
         if ({b[12],a[6]}) == loop_204[1:0]) begin
          match_flag_204 = 1'b1;
          addr[204] = loop_204[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_205 = 1'b0;
        addr[205] = 3'b0;
        for (loop_205 = 0; loop_205 < NUM_CELL; loop_205++) begin
         if ({b[13],a[6]}) == loop_205[1:0]) begin
          match_flag_205 = 1'b1;
          addr[205] = loop_205[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_206 = 1'b0;
        addr[206] = 3'b0;
        for (loop_206 = 0; loop_206 < NUM_CELL; loop_206++) begin
         if ({b[14],a[6]}) == loop_206[1:0]) begin
          match_flag_206 = 1'b1;
          addr[206] = loop_206[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_207 = 1'b0;
        addr[207] = 3'b0;
        for (loop_207 = 0; loop_207 < NUM_CELL; loop_207++) begin
         if ({b[15],a[6]}) == loop_207[1:0]) begin
          match_flag_207 = 1'b1;
          addr[207] = loop_207[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_208 = 1'b0;
        addr[208] = 3'b0;
        for (loop_208 = 0; loop_208 < NUM_CELL; loop_208++) begin
         if ({b[16],a[6]}) == loop_208[1:0]) begin
          match_flag_208 = 1'b1;
          addr[208] = loop_208[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_209 = 1'b0;
        addr[209] = 3'b0;
        for (loop_209 = 0; loop_209 < NUM_CELL; loop_209++) begin
         if ({b[17],a[6]}) == loop_209[1:0]) begin
          match_flag_209 = 1'b1;
          addr[209] = loop_209[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_210 = 1'b0;
        addr[210] = 3'b0;
        for (loop_210 = 0; loop_210 < NUM_CELL; loop_210++) begin
         if ({b[18],a[6]}) == loop_210[1:0]) begin
          match_flag_210 = 1'b1;
          addr[210] = loop_210[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_211 = 1'b0;
        addr[211] = 3'b0;
        for (loop_211 = 0; loop_211 < NUM_CELL; loop_211++) begin
         if ({b[19],a[6]}) == loop_211[1:0]) begin
          match_flag_211 = 1'b1;
          addr[211] = loop_211[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_212 = 1'b0;
        addr[212] = 3'b0;
        for (loop_212 = 0; loop_212 < NUM_CELL; loop_212++) begin
         if ({b[20],a[6]}) == loop_212[1:0]) begin
          match_flag_212 = 1'b1;
          addr[212] = loop_212[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_213 = 1'b0;
        addr[213] = 3'b0;
        for (loop_213 = 0; loop_213 < NUM_CELL; loop_213++) begin
         if ({b[21],a[6]}) == loop_213[1:0]) begin
          match_flag_213 = 1'b1;
          addr[213] = loop_213[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_214 = 1'b0;
        addr[214] = 3'b0;
        for (loop_214 = 0; loop_214 < NUM_CELL; loop_214++) begin
         if ({b[22],a[6]}) == loop_214[1:0]) begin
          match_flag_214 = 1'b1;
          addr[214] = loop_214[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_215 = 1'b0;
        addr[215] = 3'b0;
        for (loop_215 = 0; loop_215 < NUM_CELL; loop_215++) begin
         if ({b[23],a[6]}) == loop_215[1:0]) begin
          match_flag_215 = 1'b1;
          addr[215] = loop_215[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_216 = 1'b0;
        addr[216] = 3'b0;
        for (loop_216 = 0; loop_216 < NUM_CELL; loop_216++) begin
         if ({b[24],a[6]}) == loop_216[1:0]) begin
          match_flag_216 = 1'b1;
          addr[216] = loop_216[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_217 = 1'b0;
        addr[217] = 3'b0;
        for (loop_217 = 0; loop_217 < NUM_CELL; loop_217++) begin
         if ({b[25],a[6]}) == loop_217[1:0]) begin
          match_flag_217 = 1'b1;
          addr[217] = loop_217[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_218 = 1'b0;
        addr[218] = 3'b0;
        for (loop_218 = 0; loop_218 < NUM_CELL; loop_218++) begin
         if ({b[26],a[6]}) == loop_218[1:0]) begin
          match_flag_218 = 1'b1;
          addr[218] = loop_218[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_219 = 1'b0;
        addr[219] = 3'b0;
        for (loop_219 = 0; loop_219 < NUM_CELL; loop_219++) begin
         if ({b[27],a[6]}) == loop_219[1:0]) begin
          match_flag_219 = 1'b1;
          addr[219] = loop_219[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_220 = 1'b0;
        addr[220] = 3'b0;
        for (loop_220 = 0; loop_220 < NUM_CELL; loop_220++) begin
         if ({b[28],a[6]}) == loop_220[1:0]) begin
          match_flag_220 = 1'b1;
          addr[220] = loop_220[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_221 = 1'b0;
        addr[221] = 3'b0;
        for (loop_221 = 0; loop_221 < NUM_CELL; loop_221++) begin
         if ({b[29],a[6]}) == loop_221[1:0]) begin
          match_flag_221 = 1'b1;
          addr[221] = loop_221[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_222 = 1'b0;
        addr[222] = 3'b0;
        for (loop_222 = 0; loop_222 < NUM_CELL; loop_222++) begin
         if ({b[30],a[6]}) == loop_222[1:0]) begin
          match_flag_222 = 1'b1;
          addr[222] = loop_222[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_223 = 1'b0;
        addr[223] = 3'b0;
        for (loop_223 = 0; loop_223 < NUM_CELL; loop_223++) begin
         if ({b[31],a[6]}) == loop_223[1:0]) begin
          match_flag_223 = 1'b1;
          addr[223] = loop_223[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_224 = 1'b0;
        addr[224] = 3'b0;
        for (loop_224 = 0; loop_224 < NUM_CELL; loop_224++) begin
         if ({b[0],a[7]}) == loop_224[1:0]) begin
          match_flag_224 = 1'b1;
          addr[224] = loop_224[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_225 = 1'b0;
        addr[225] = 3'b0;
        for (loop_225 = 0; loop_225 < NUM_CELL; loop_225++) begin
         if ({b[1],a[7]}) == loop_225[1:0]) begin
          match_flag_225 = 1'b1;
          addr[225] = loop_225[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_226 = 1'b0;
        addr[226] = 3'b0;
        for (loop_226 = 0; loop_226 < NUM_CELL; loop_226++) begin
         if ({b[2],a[7]}) == loop_226[1:0]) begin
          match_flag_226 = 1'b1;
          addr[226] = loop_226[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_227 = 1'b0;
        addr[227] = 3'b0;
        for (loop_227 = 0; loop_227 < NUM_CELL; loop_227++) begin
         if ({b[3],a[7]}) == loop_227[1:0]) begin
          match_flag_227 = 1'b1;
          addr[227] = loop_227[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_228 = 1'b0;
        addr[228] = 3'b0;
        for (loop_228 = 0; loop_228 < NUM_CELL; loop_228++) begin
         if ({b[4],a[7]}) == loop_228[1:0]) begin
          match_flag_228 = 1'b1;
          addr[228] = loop_228[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_229 = 1'b0;
        addr[229] = 3'b0;
        for (loop_229 = 0; loop_229 < NUM_CELL; loop_229++) begin
         if ({b[5],a[7]}) == loop_229[1:0]) begin
          match_flag_229 = 1'b1;
          addr[229] = loop_229[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_230 = 1'b0;
        addr[230] = 3'b0;
        for (loop_230 = 0; loop_230 < NUM_CELL; loop_230++) begin
         if ({b[6],a[7]}) == loop_230[1:0]) begin
          match_flag_230 = 1'b1;
          addr[230] = loop_230[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_231 = 1'b0;
        addr[231] = 3'b0;
        for (loop_231 = 0; loop_231 < NUM_CELL; loop_231++) begin
         if ({b[7],a[7]}) == loop_231[1:0]) begin
          match_flag_231 = 1'b1;
          addr[231] = loop_231[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_232 = 1'b0;
        addr[232] = 3'b0;
        for (loop_232 = 0; loop_232 < NUM_CELL; loop_232++) begin
         if ({b[8],a[7]}) == loop_232[1:0]) begin
          match_flag_232 = 1'b1;
          addr[232] = loop_232[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_233 = 1'b0;
        addr[233] = 3'b0;
        for (loop_233 = 0; loop_233 < NUM_CELL; loop_233++) begin
         if ({b[9],a[7]}) == loop_233[1:0]) begin
          match_flag_233 = 1'b1;
          addr[233] = loop_233[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_234 = 1'b0;
        addr[234] = 3'b0;
        for (loop_234 = 0; loop_234 < NUM_CELL; loop_234++) begin
         if ({b[10],a[7]}) == loop_234[1:0]) begin
          match_flag_234 = 1'b1;
          addr[234] = loop_234[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_235 = 1'b0;
        addr[235] = 3'b0;
        for (loop_235 = 0; loop_235 < NUM_CELL; loop_235++) begin
         if ({b[11],a[7]}) == loop_235[1:0]) begin
          match_flag_235 = 1'b1;
          addr[235] = loop_235[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_236 = 1'b0;
        addr[236] = 3'b0;
        for (loop_236 = 0; loop_236 < NUM_CELL; loop_236++) begin
         if ({b[12],a[7]}) == loop_236[1:0]) begin
          match_flag_236 = 1'b1;
          addr[236] = loop_236[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_237 = 1'b0;
        addr[237] = 3'b0;
        for (loop_237 = 0; loop_237 < NUM_CELL; loop_237++) begin
         if ({b[13],a[7]}) == loop_237[1:0]) begin
          match_flag_237 = 1'b1;
          addr[237] = loop_237[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_238 = 1'b0;
        addr[238] = 3'b0;
        for (loop_238 = 0; loop_238 < NUM_CELL; loop_238++) begin
         if ({b[14],a[7]}) == loop_238[1:0]) begin
          match_flag_238 = 1'b1;
          addr[238] = loop_238[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_239 = 1'b0;
        addr[239] = 3'b0;
        for (loop_239 = 0; loop_239 < NUM_CELL; loop_239++) begin
         if ({b[15],a[7]}) == loop_239[1:0]) begin
          match_flag_239 = 1'b1;
          addr[239] = loop_239[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_240 = 1'b0;
        addr[240] = 3'b0;
        for (loop_240 = 0; loop_240 < NUM_CELL; loop_240++) begin
         if ({b[16],a[7]}) == loop_240[1:0]) begin
          match_flag_240 = 1'b1;
          addr[240] = loop_240[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_241 = 1'b0;
        addr[241] = 3'b0;
        for (loop_241 = 0; loop_241 < NUM_CELL; loop_241++) begin
         if ({b[17],a[7]}) == loop_241[1:0]) begin
          match_flag_241 = 1'b1;
          addr[241] = loop_241[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_242 = 1'b0;
        addr[242] = 3'b0;
        for (loop_242 = 0; loop_242 < NUM_CELL; loop_242++) begin
         if ({b[18],a[7]}) == loop_242[1:0]) begin
          match_flag_242 = 1'b1;
          addr[242] = loop_242[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_243 = 1'b0;
        addr[243] = 3'b0;
        for (loop_243 = 0; loop_243 < NUM_CELL; loop_243++) begin
         if ({b[19],a[7]}) == loop_243[1:0]) begin
          match_flag_243 = 1'b1;
          addr[243] = loop_243[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_244 = 1'b0;
        addr[244] = 3'b0;
        for (loop_244 = 0; loop_244 < NUM_CELL; loop_244++) begin
         if ({b[20],a[7]}) == loop_244[1:0]) begin
          match_flag_244 = 1'b1;
          addr[244] = loop_244[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_245 = 1'b0;
        addr[245] = 3'b0;
        for (loop_245 = 0; loop_245 < NUM_CELL; loop_245++) begin
         if ({b[21],a[7]}) == loop_245[1:0]) begin
          match_flag_245 = 1'b1;
          addr[245] = loop_245[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_246 = 1'b0;
        addr[246] = 3'b0;
        for (loop_246 = 0; loop_246 < NUM_CELL; loop_246++) begin
         if ({b[22],a[7]}) == loop_246[1:0]) begin
          match_flag_246 = 1'b1;
          addr[246] = loop_246[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_247 = 1'b0;
        addr[247] = 3'b0;
        for (loop_247 = 0; loop_247 < NUM_CELL; loop_247++) begin
         if ({b[23],a[7]}) == loop_247[1:0]) begin
          match_flag_247 = 1'b1;
          addr[247] = loop_247[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_248 = 1'b0;
        addr[248] = 3'b0;
        for (loop_248 = 0; loop_248 < NUM_CELL; loop_248++) begin
         if ({b[24],a[7]}) == loop_248[1:0]) begin
          match_flag_248 = 1'b1;
          addr[248] = loop_248[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_249 = 1'b0;
        addr[249] = 3'b0;
        for (loop_249 = 0; loop_249 < NUM_CELL; loop_249++) begin
         if ({b[25],a[7]}) == loop_249[1:0]) begin
          match_flag_249 = 1'b1;
          addr[249] = loop_249[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_250 = 1'b0;
        addr[250] = 3'b0;
        for (loop_250 = 0; loop_250 < NUM_CELL; loop_250++) begin
         if ({b[26],a[7]}) == loop_250[1:0]) begin
          match_flag_250 = 1'b1;
          addr[250] = loop_250[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_251 = 1'b0;
        addr[251] = 3'b0;
        for (loop_251 = 0; loop_251 < NUM_CELL; loop_251++) begin
         if ({b[27],a[7]}) == loop_251[1:0]) begin
          match_flag_251 = 1'b1;
          addr[251] = loop_251[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_252 = 1'b0;
        addr[252] = 3'b0;
        for (loop_252 = 0; loop_252 < NUM_CELL; loop_252++) begin
         if ({b[28],a[7]}) == loop_252[1:0]) begin
          match_flag_252 = 1'b1;
          addr[252] = loop_252[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_253 = 1'b0;
        addr[253] = 3'b0;
        for (loop_253 = 0; loop_253 < NUM_CELL; loop_253++) begin
         if ({b[29],a[7]}) == loop_253[1:0]) begin
          match_flag_253 = 1'b1;
          addr[253] = loop_253[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_254 = 1'b0;
        addr[254] = 3'b0;
        for (loop_254 = 0; loop_254 < NUM_CELL; loop_254++) begin
         if ({b[30],a[7]}) == loop_254[1:0]) begin
          match_flag_254 = 1'b1;
          addr[254] = loop_254[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_255 = 1'b0;
        addr[255] = 3'b0;
        for (loop_255 = 0; loop_255 < NUM_CELL; loop_255++) begin
         if ({b[31],a[7]}) == loop_255[1:0]) begin
          match_flag_255 = 1'b1;
          addr[255] = loop_255[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_256 = 1'b0;
        addr[256] = 3'b0;
        for (loop_256 = 0; loop_256 < NUM_CELL; loop_256++) begin
         if ({b[0],a[8]}) == loop_256[1:0]) begin
          match_flag_256 = 1'b1;
          addr[256] = loop_256[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_257 = 1'b0;
        addr[257] = 3'b0;
        for (loop_257 = 0; loop_257 < NUM_CELL; loop_257++) begin
         if ({b[1],a[8]}) == loop_257[1:0]) begin
          match_flag_257 = 1'b1;
          addr[257] = loop_257[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_258 = 1'b0;
        addr[258] = 3'b0;
        for (loop_258 = 0; loop_258 < NUM_CELL; loop_258++) begin
         if ({b[2],a[8]}) == loop_258[1:0]) begin
          match_flag_258 = 1'b1;
          addr[258] = loop_258[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_259 = 1'b0;
        addr[259] = 3'b0;
        for (loop_259 = 0; loop_259 < NUM_CELL; loop_259++) begin
         if ({b[3],a[8]}) == loop_259[1:0]) begin
          match_flag_259 = 1'b1;
          addr[259] = loop_259[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_260 = 1'b0;
        addr[260] = 3'b0;
        for (loop_260 = 0; loop_260 < NUM_CELL; loop_260++) begin
         if ({b[4],a[8]}) == loop_260[1:0]) begin
          match_flag_260 = 1'b1;
          addr[260] = loop_260[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_261 = 1'b0;
        addr[261] = 3'b0;
        for (loop_261 = 0; loop_261 < NUM_CELL; loop_261++) begin
         if ({b[5],a[8]}) == loop_261[1:0]) begin
          match_flag_261 = 1'b1;
          addr[261] = loop_261[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_262 = 1'b0;
        addr[262] = 3'b0;
        for (loop_262 = 0; loop_262 < NUM_CELL; loop_262++) begin
         if ({b[6],a[8]}) == loop_262[1:0]) begin
          match_flag_262 = 1'b1;
          addr[262] = loop_262[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_263 = 1'b0;
        addr[263] = 3'b0;
        for (loop_263 = 0; loop_263 < NUM_CELL; loop_263++) begin
         if ({b[7],a[8]}) == loop_263[1:0]) begin
          match_flag_263 = 1'b1;
          addr[263] = loop_263[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_264 = 1'b0;
        addr[264] = 3'b0;
        for (loop_264 = 0; loop_264 < NUM_CELL; loop_264++) begin
         if ({b[8],a[8]}) == loop_264[1:0]) begin
          match_flag_264 = 1'b1;
          addr[264] = loop_264[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_265 = 1'b0;
        addr[265] = 3'b0;
        for (loop_265 = 0; loop_265 < NUM_CELL; loop_265++) begin
         if ({b[9],a[8]}) == loop_265[1:0]) begin
          match_flag_265 = 1'b1;
          addr[265] = loop_265[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_266 = 1'b0;
        addr[266] = 3'b0;
        for (loop_266 = 0; loop_266 < NUM_CELL; loop_266++) begin
         if ({b[10],a[8]}) == loop_266[1:0]) begin
          match_flag_266 = 1'b1;
          addr[266] = loop_266[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_267 = 1'b0;
        addr[267] = 3'b0;
        for (loop_267 = 0; loop_267 < NUM_CELL; loop_267++) begin
         if ({b[11],a[8]}) == loop_267[1:0]) begin
          match_flag_267 = 1'b1;
          addr[267] = loop_267[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_268 = 1'b0;
        addr[268] = 3'b0;
        for (loop_268 = 0; loop_268 < NUM_CELL; loop_268++) begin
         if ({b[12],a[8]}) == loop_268[1:0]) begin
          match_flag_268 = 1'b1;
          addr[268] = loop_268[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_269 = 1'b0;
        addr[269] = 3'b0;
        for (loop_269 = 0; loop_269 < NUM_CELL; loop_269++) begin
         if ({b[13],a[8]}) == loop_269[1:0]) begin
          match_flag_269 = 1'b1;
          addr[269] = loop_269[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_270 = 1'b0;
        addr[270] = 3'b0;
        for (loop_270 = 0; loop_270 < NUM_CELL; loop_270++) begin
         if ({b[14],a[8]}) == loop_270[1:0]) begin
          match_flag_270 = 1'b1;
          addr[270] = loop_270[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_271 = 1'b0;
        addr[271] = 3'b0;
        for (loop_271 = 0; loop_271 < NUM_CELL; loop_271++) begin
         if ({b[15],a[8]}) == loop_271[1:0]) begin
          match_flag_271 = 1'b1;
          addr[271] = loop_271[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_272 = 1'b0;
        addr[272] = 3'b0;
        for (loop_272 = 0; loop_272 < NUM_CELL; loop_272++) begin
         if ({b[16],a[8]}) == loop_272[1:0]) begin
          match_flag_272 = 1'b1;
          addr[272] = loop_272[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_273 = 1'b0;
        addr[273] = 3'b0;
        for (loop_273 = 0; loop_273 < NUM_CELL; loop_273++) begin
         if ({b[17],a[8]}) == loop_273[1:0]) begin
          match_flag_273 = 1'b1;
          addr[273] = loop_273[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_274 = 1'b0;
        addr[274] = 3'b0;
        for (loop_274 = 0; loop_274 < NUM_CELL; loop_274++) begin
         if ({b[18],a[8]}) == loop_274[1:0]) begin
          match_flag_274 = 1'b1;
          addr[274] = loop_274[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_275 = 1'b0;
        addr[275] = 3'b0;
        for (loop_275 = 0; loop_275 < NUM_CELL; loop_275++) begin
         if ({b[19],a[8]}) == loop_275[1:0]) begin
          match_flag_275 = 1'b1;
          addr[275] = loop_275[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_276 = 1'b0;
        addr[276] = 3'b0;
        for (loop_276 = 0; loop_276 < NUM_CELL; loop_276++) begin
         if ({b[20],a[8]}) == loop_276[1:0]) begin
          match_flag_276 = 1'b1;
          addr[276] = loop_276[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_277 = 1'b0;
        addr[277] = 3'b0;
        for (loop_277 = 0; loop_277 < NUM_CELL; loop_277++) begin
         if ({b[21],a[8]}) == loop_277[1:0]) begin
          match_flag_277 = 1'b1;
          addr[277] = loop_277[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_278 = 1'b0;
        addr[278] = 3'b0;
        for (loop_278 = 0; loop_278 < NUM_CELL; loop_278++) begin
         if ({b[22],a[8]}) == loop_278[1:0]) begin
          match_flag_278 = 1'b1;
          addr[278] = loop_278[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_279 = 1'b0;
        addr[279] = 3'b0;
        for (loop_279 = 0; loop_279 < NUM_CELL; loop_279++) begin
         if ({b[23],a[8]}) == loop_279[1:0]) begin
          match_flag_279 = 1'b1;
          addr[279] = loop_279[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_280 = 1'b0;
        addr[280] = 3'b0;
        for (loop_280 = 0; loop_280 < NUM_CELL; loop_280++) begin
         if ({b[24],a[8]}) == loop_280[1:0]) begin
          match_flag_280 = 1'b1;
          addr[280] = loop_280[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_281 = 1'b0;
        addr[281] = 3'b0;
        for (loop_281 = 0; loop_281 < NUM_CELL; loop_281++) begin
         if ({b[25],a[8]}) == loop_281[1:0]) begin
          match_flag_281 = 1'b1;
          addr[281] = loop_281[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_282 = 1'b0;
        addr[282] = 3'b0;
        for (loop_282 = 0; loop_282 < NUM_CELL; loop_282++) begin
         if ({b[26],a[8]}) == loop_282[1:0]) begin
          match_flag_282 = 1'b1;
          addr[282] = loop_282[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_283 = 1'b0;
        addr[283] = 3'b0;
        for (loop_283 = 0; loop_283 < NUM_CELL; loop_283++) begin
         if ({b[27],a[8]}) == loop_283[1:0]) begin
          match_flag_283 = 1'b1;
          addr[283] = loop_283[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_284 = 1'b0;
        addr[284] = 3'b0;
        for (loop_284 = 0; loop_284 < NUM_CELL; loop_284++) begin
         if ({b[28],a[8]}) == loop_284[1:0]) begin
          match_flag_284 = 1'b1;
          addr[284] = loop_284[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_285 = 1'b0;
        addr[285] = 3'b0;
        for (loop_285 = 0; loop_285 < NUM_CELL; loop_285++) begin
         if ({b[29],a[8]}) == loop_285[1:0]) begin
          match_flag_285 = 1'b1;
          addr[285] = loop_285[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_286 = 1'b0;
        addr[286] = 3'b0;
        for (loop_286 = 0; loop_286 < NUM_CELL; loop_286++) begin
         if ({b[30],a[8]}) == loop_286[1:0]) begin
          match_flag_286 = 1'b1;
          addr[286] = loop_286[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_287 = 1'b0;
        addr[287] = 3'b0;
        for (loop_287 = 0; loop_287 < NUM_CELL; loop_287++) begin
         if ({b[31],a[8]}) == loop_287[1:0]) begin
          match_flag_287 = 1'b1;
          addr[287] = loop_287[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_288 = 1'b0;
        addr[288] = 3'b0;
        for (loop_288 = 0; loop_288 < NUM_CELL; loop_288++) begin
         if ({b[0],a[9]}) == loop_288[1:0]) begin
          match_flag_288 = 1'b1;
          addr[288] = loop_288[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_289 = 1'b0;
        addr[289] = 3'b0;
        for (loop_289 = 0; loop_289 < NUM_CELL; loop_289++) begin
         if ({b[1],a[9]}) == loop_289[1:0]) begin
          match_flag_289 = 1'b1;
          addr[289] = loop_289[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_290 = 1'b0;
        addr[290] = 3'b0;
        for (loop_290 = 0; loop_290 < NUM_CELL; loop_290++) begin
         if ({b[2],a[9]}) == loop_290[1:0]) begin
          match_flag_290 = 1'b1;
          addr[290] = loop_290[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_291 = 1'b0;
        addr[291] = 3'b0;
        for (loop_291 = 0; loop_291 < NUM_CELL; loop_291++) begin
         if ({b[3],a[9]}) == loop_291[1:0]) begin
          match_flag_291 = 1'b1;
          addr[291] = loop_291[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_292 = 1'b0;
        addr[292] = 3'b0;
        for (loop_292 = 0; loop_292 < NUM_CELL; loop_292++) begin
         if ({b[4],a[9]}) == loop_292[1:0]) begin
          match_flag_292 = 1'b1;
          addr[292] = loop_292[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_293 = 1'b0;
        addr[293] = 3'b0;
        for (loop_293 = 0; loop_293 < NUM_CELL; loop_293++) begin
         if ({b[5],a[9]}) == loop_293[1:0]) begin
          match_flag_293 = 1'b1;
          addr[293] = loop_293[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_294 = 1'b0;
        addr[294] = 3'b0;
        for (loop_294 = 0; loop_294 < NUM_CELL; loop_294++) begin
         if ({b[6],a[9]}) == loop_294[1:0]) begin
          match_flag_294 = 1'b1;
          addr[294] = loop_294[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_295 = 1'b0;
        addr[295] = 3'b0;
        for (loop_295 = 0; loop_295 < NUM_CELL; loop_295++) begin
         if ({b[7],a[9]}) == loop_295[1:0]) begin
          match_flag_295 = 1'b1;
          addr[295] = loop_295[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_296 = 1'b0;
        addr[296] = 3'b0;
        for (loop_296 = 0; loop_296 < NUM_CELL; loop_296++) begin
         if ({b[8],a[9]}) == loop_296[1:0]) begin
          match_flag_296 = 1'b1;
          addr[296] = loop_296[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_297 = 1'b0;
        addr[297] = 3'b0;
        for (loop_297 = 0; loop_297 < NUM_CELL; loop_297++) begin
         if ({b[9],a[9]}) == loop_297[1:0]) begin
          match_flag_297 = 1'b1;
          addr[297] = loop_297[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_298 = 1'b0;
        addr[298] = 3'b0;
        for (loop_298 = 0; loop_298 < NUM_CELL; loop_298++) begin
         if ({b[10],a[9]}) == loop_298[1:0]) begin
          match_flag_298 = 1'b1;
          addr[298] = loop_298[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_299 = 1'b0;
        addr[299] = 3'b0;
        for (loop_299 = 0; loop_299 < NUM_CELL; loop_299++) begin
         if ({b[11],a[9]}) == loop_299[1:0]) begin
          match_flag_299 = 1'b1;
          addr[299] = loop_299[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_300 = 1'b0;
        addr[300] = 3'b0;
        for (loop_300 = 0; loop_300 < NUM_CELL; loop_300++) begin
         if ({b[12],a[9]}) == loop_300[1:0]) begin
          match_flag_300 = 1'b1;
          addr[300] = loop_300[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_301 = 1'b0;
        addr[301] = 3'b0;
        for (loop_301 = 0; loop_301 < NUM_CELL; loop_301++) begin
         if ({b[13],a[9]}) == loop_301[1:0]) begin
          match_flag_301 = 1'b1;
          addr[301] = loop_301[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_302 = 1'b0;
        addr[302] = 3'b0;
        for (loop_302 = 0; loop_302 < NUM_CELL; loop_302++) begin
         if ({b[14],a[9]}) == loop_302[1:0]) begin
          match_flag_302 = 1'b1;
          addr[302] = loop_302[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_303 = 1'b0;
        addr[303] = 3'b0;
        for (loop_303 = 0; loop_303 < NUM_CELL; loop_303++) begin
         if ({b[15],a[9]}) == loop_303[1:0]) begin
          match_flag_303 = 1'b1;
          addr[303] = loop_303[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_304 = 1'b0;
        addr[304] = 3'b0;
        for (loop_304 = 0; loop_304 < NUM_CELL; loop_304++) begin
         if ({b[16],a[9]}) == loop_304[1:0]) begin
          match_flag_304 = 1'b1;
          addr[304] = loop_304[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_305 = 1'b0;
        addr[305] = 3'b0;
        for (loop_305 = 0; loop_305 < NUM_CELL; loop_305++) begin
         if ({b[17],a[9]}) == loop_305[1:0]) begin
          match_flag_305 = 1'b1;
          addr[305] = loop_305[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_306 = 1'b0;
        addr[306] = 3'b0;
        for (loop_306 = 0; loop_306 < NUM_CELL; loop_306++) begin
         if ({b[18],a[9]}) == loop_306[1:0]) begin
          match_flag_306 = 1'b1;
          addr[306] = loop_306[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_307 = 1'b0;
        addr[307] = 3'b0;
        for (loop_307 = 0; loop_307 < NUM_CELL; loop_307++) begin
         if ({b[19],a[9]}) == loop_307[1:0]) begin
          match_flag_307 = 1'b1;
          addr[307] = loop_307[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_308 = 1'b0;
        addr[308] = 3'b0;
        for (loop_308 = 0; loop_308 < NUM_CELL; loop_308++) begin
         if ({b[20],a[9]}) == loop_308[1:0]) begin
          match_flag_308 = 1'b1;
          addr[308] = loop_308[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_309 = 1'b0;
        addr[309] = 3'b0;
        for (loop_309 = 0; loop_309 < NUM_CELL; loop_309++) begin
         if ({b[21],a[9]}) == loop_309[1:0]) begin
          match_flag_309 = 1'b1;
          addr[309] = loop_309[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_310 = 1'b0;
        addr[310] = 3'b0;
        for (loop_310 = 0; loop_310 < NUM_CELL; loop_310++) begin
         if ({b[22],a[9]}) == loop_310[1:0]) begin
          match_flag_310 = 1'b1;
          addr[310] = loop_310[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_311 = 1'b0;
        addr[311] = 3'b0;
        for (loop_311 = 0; loop_311 < NUM_CELL; loop_311++) begin
         if ({b[23],a[9]}) == loop_311[1:0]) begin
          match_flag_311 = 1'b1;
          addr[311] = loop_311[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_312 = 1'b0;
        addr[312] = 3'b0;
        for (loop_312 = 0; loop_312 < NUM_CELL; loop_312++) begin
         if ({b[24],a[9]}) == loop_312[1:0]) begin
          match_flag_312 = 1'b1;
          addr[312] = loop_312[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_313 = 1'b0;
        addr[313] = 3'b0;
        for (loop_313 = 0; loop_313 < NUM_CELL; loop_313++) begin
         if ({b[25],a[9]}) == loop_313[1:0]) begin
          match_flag_313 = 1'b1;
          addr[313] = loop_313[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_314 = 1'b0;
        addr[314] = 3'b0;
        for (loop_314 = 0; loop_314 < NUM_CELL; loop_314++) begin
         if ({b[26],a[9]}) == loop_314[1:0]) begin
          match_flag_314 = 1'b1;
          addr[314] = loop_314[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_315 = 1'b0;
        addr[315] = 3'b0;
        for (loop_315 = 0; loop_315 < NUM_CELL; loop_315++) begin
         if ({b[27],a[9]}) == loop_315[1:0]) begin
          match_flag_315 = 1'b1;
          addr[315] = loop_315[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_316 = 1'b0;
        addr[316] = 3'b0;
        for (loop_316 = 0; loop_316 < NUM_CELL; loop_316++) begin
         if ({b[28],a[9]}) == loop_316[1:0]) begin
          match_flag_316 = 1'b1;
          addr[316] = loop_316[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_317 = 1'b0;
        addr[317] = 3'b0;
        for (loop_317 = 0; loop_317 < NUM_CELL; loop_317++) begin
         if ({b[29],a[9]}) == loop_317[1:0]) begin
          match_flag_317 = 1'b1;
          addr[317] = loop_317[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_318 = 1'b0;
        addr[318] = 3'b0;
        for (loop_318 = 0; loop_318 < NUM_CELL; loop_318++) begin
         if ({b[30],a[9]}) == loop_318[1:0]) begin
          match_flag_318 = 1'b1;
          addr[318] = loop_318[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_319 = 1'b0;
        addr[319] = 3'b0;
        for (loop_319 = 0; loop_319 < NUM_CELL; loop_319++) begin
         if ({b[31],a[9]}) == loop_319[1:0]) begin
          match_flag_319 = 1'b1;
          addr[319] = loop_319[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_320 = 1'b0;
        addr[320] = 3'b0;
        for (loop_320 = 0; loop_320 < NUM_CELL; loop_320++) begin
         if ({b[0],a[10]}) == loop_320[1:0]) begin
          match_flag_320 = 1'b1;
          addr[320] = loop_320[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_321 = 1'b0;
        addr[321] = 3'b0;
        for (loop_321 = 0; loop_321 < NUM_CELL; loop_321++) begin
         if ({b[1],a[10]}) == loop_321[1:0]) begin
          match_flag_321 = 1'b1;
          addr[321] = loop_321[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_322 = 1'b0;
        addr[322] = 3'b0;
        for (loop_322 = 0; loop_322 < NUM_CELL; loop_322++) begin
         if ({b[2],a[10]}) == loop_322[1:0]) begin
          match_flag_322 = 1'b1;
          addr[322] = loop_322[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_323 = 1'b0;
        addr[323] = 3'b0;
        for (loop_323 = 0; loop_323 < NUM_CELL; loop_323++) begin
         if ({b[3],a[10]}) == loop_323[1:0]) begin
          match_flag_323 = 1'b1;
          addr[323] = loop_323[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_324 = 1'b0;
        addr[324] = 3'b0;
        for (loop_324 = 0; loop_324 < NUM_CELL; loop_324++) begin
         if ({b[4],a[10]}) == loop_324[1:0]) begin
          match_flag_324 = 1'b1;
          addr[324] = loop_324[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_325 = 1'b0;
        addr[325] = 3'b0;
        for (loop_325 = 0; loop_325 < NUM_CELL; loop_325++) begin
         if ({b[5],a[10]}) == loop_325[1:0]) begin
          match_flag_325 = 1'b1;
          addr[325] = loop_325[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_326 = 1'b0;
        addr[326] = 3'b0;
        for (loop_326 = 0; loop_326 < NUM_CELL; loop_326++) begin
         if ({b[6],a[10]}) == loop_326[1:0]) begin
          match_flag_326 = 1'b1;
          addr[326] = loop_326[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_327 = 1'b0;
        addr[327] = 3'b0;
        for (loop_327 = 0; loop_327 < NUM_CELL; loop_327++) begin
         if ({b[7],a[10]}) == loop_327[1:0]) begin
          match_flag_327 = 1'b1;
          addr[327] = loop_327[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_328 = 1'b0;
        addr[328] = 3'b0;
        for (loop_328 = 0; loop_328 < NUM_CELL; loop_328++) begin
         if ({b[8],a[10]}) == loop_328[1:0]) begin
          match_flag_328 = 1'b1;
          addr[328] = loop_328[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_329 = 1'b0;
        addr[329] = 3'b0;
        for (loop_329 = 0; loop_329 < NUM_CELL; loop_329++) begin
         if ({b[9],a[10]}) == loop_329[1:0]) begin
          match_flag_329 = 1'b1;
          addr[329] = loop_329[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_330 = 1'b0;
        addr[330] = 3'b0;
        for (loop_330 = 0; loop_330 < NUM_CELL; loop_330++) begin
         if ({b[10],a[10]}) == loop_330[1:0]) begin
          match_flag_330 = 1'b1;
          addr[330] = loop_330[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_331 = 1'b0;
        addr[331] = 3'b0;
        for (loop_331 = 0; loop_331 < NUM_CELL; loop_331++) begin
         if ({b[11],a[10]}) == loop_331[1:0]) begin
          match_flag_331 = 1'b1;
          addr[331] = loop_331[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_332 = 1'b0;
        addr[332] = 3'b0;
        for (loop_332 = 0; loop_332 < NUM_CELL; loop_332++) begin
         if ({b[12],a[10]}) == loop_332[1:0]) begin
          match_flag_332 = 1'b1;
          addr[332] = loop_332[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_333 = 1'b0;
        addr[333] = 3'b0;
        for (loop_333 = 0; loop_333 < NUM_CELL; loop_333++) begin
         if ({b[13],a[10]}) == loop_333[1:0]) begin
          match_flag_333 = 1'b1;
          addr[333] = loop_333[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_334 = 1'b0;
        addr[334] = 3'b0;
        for (loop_334 = 0; loop_334 < NUM_CELL; loop_334++) begin
         if ({b[14],a[10]}) == loop_334[1:0]) begin
          match_flag_334 = 1'b1;
          addr[334] = loop_334[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_335 = 1'b0;
        addr[335] = 3'b0;
        for (loop_335 = 0; loop_335 < NUM_CELL; loop_335++) begin
         if ({b[15],a[10]}) == loop_335[1:0]) begin
          match_flag_335 = 1'b1;
          addr[335] = loop_335[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_336 = 1'b0;
        addr[336] = 3'b0;
        for (loop_336 = 0; loop_336 < NUM_CELL; loop_336++) begin
         if ({b[16],a[10]}) == loop_336[1:0]) begin
          match_flag_336 = 1'b1;
          addr[336] = loop_336[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_337 = 1'b0;
        addr[337] = 3'b0;
        for (loop_337 = 0; loop_337 < NUM_CELL; loop_337++) begin
         if ({b[17],a[10]}) == loop_337[1:0]) begin
          match_flag_337 = 1'b1;
          addr[337] = loop_337[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_338 = 1'b0;
        addr[338] = 3'b0;
        for (loop_338 = 0; loop_338 < NUM_CELL; loop_338++) begin
         if ({b[18],a[10]}) == loop_338[1:0]) begin
          match_flag_338 = 1'b1;
          addr[338] = loop_338[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_339 = 1'b0;
        addr[339] = 3'b0;
        for (loop_339 = 0; loop_339 < NUM_CELL; loop_339++) begin
         if ({b[19],a[10]}) == loop_339[1:0]) begin
          match_flag_339 = 1'b1;
          addr[339] = loop_339[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_340 = 1'b0;
        addr[340] = 3'b0;
        for (loop_340 = 0; loop_340 < NUM_CELL; loop_340++) begin
         if ({b[20],a[10]}) == loop_340[1:0]) begin
          match_flag_340 = 1'b1;
          addr[340] = loop_340[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_341 = 1'b0;
        addr[341] = 3'b0;
        for (loop_341 = 0; loop_341 < NUM_CELL; loop_341++) begin
         if ({b[21],a[10]}) == loop_341[1:0]) begin
          match_flag_341 = 1'b1;
          addr[341] = loop_341[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_342 = 1'b0;
        addr[342] = 3'b0;
        for (loop_342 = 0; loop_342 < NUM_CELL; loop_342++) begin
         if ({b[22],a[10]}) == loop_342[1:0]) begin
          match_flag_342 = 1'b1;
          addr[342] = loop_342[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_343 = 1'b0;
        addr[343] = 3'b0;
        for (loop_343 = 0; loop_343 < NUM_CELL; loop_343++) begin
         if ({b[23],a[10]}) == loop_343[1:0]) begin
          match_flag_343 = 1'b1;
          addr[343] = loop_343[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_344 = 1'b0;
        addr[344] = 3'b0;
        for (loop_344 = 0; loop_344 < NUM_CELL; loop_344++) begin
         if ({b[24],a[10]}) == loop_344[1:0]) begin
          match_flag_344 = 1'b1;
          addr[344] = loop_344[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_345 = 1'b0;
        addr[345] = 3'b0;
        for (loop_345 = 0; loop_345 < NUM_CELL; loop_345++) begin
         if ({b[25],a[10]}) == loop_345[1:0]) begin
          match_flag_345 = 1'b1;
          addr[345] = loop_345[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_346 = 1'b0;
        addr[346] = 3'b0;
        for (loop_346 = 0; loop_346 < NUM_CELL; loop_346++) begin
         if ({b[26],a[10]}) == loop_346[1:0]) begin
          match_flag_346 = 1'b1;
          addr[346] = loop_346[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_347 = 1'b0;
        addr[347] = 3'b0;
        for (loop_347 = 0; loop_347 < NUM_CELL; loop_347++) begin
         if ({b[27],a[10]}) == loop_347[1:0]) begin
          match_flag_347 = 1'b1;
          addr[347] = loop_347[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_348 = 1'b0;
        addr[348] = 3'b0;
        for (loop_348 = 0; loop_348 < NUM_CELL; loop_348++) begin
         if ({b[28],a[10]}) == loop_348[1:0]) begin
          match_flag_348 = 1'b1;
          addr[348] = loop_348[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_349 = 1'b0;
        addr[349] = 3'b0;
        for (loop_349 = 0; loop_349 < NUM_CELL; loop_349++) begin
         if ({b[29],a[10]}) == loop_349[1:0]) begin
          match_flag_349 = 1'b1;
          addr[349] = loop_349[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_350 = 1'b0;
        addr[350] = 3'b0;
        for (loop_350 = 0; loop_350 < NUM_CELL; loop_350++) begin
         if ({b[30],a[10]}) == loop_350[1:0]) begin
          match_flag_350 = 1'b1;
          addr[350] = loop_350[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_351 = 1'b0;
        addr[351] = 3'b0;
        for (loop_351 = 0; loop_351 < NUM_CELL; loop_351++) begin
         if ({b[31],a[10]}) == loop_351[1:0]) begin
          match_flag_351 = 1'b1;
          addr[351] = loop_351[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_352 = 1'b0;
        addr[352] = 3'b0;
        for (loop_352 = 0; loop_352 < NUM_CELL; loop_352++) begin
         if ({b[0],a[11]}) == loop_352[1:0]) begin
          match_flag_352 = 1'b1;
          addr[352] = loop_352[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_353 = 1'b0;
        addr[353] = 3'b0;
        for (loop_353 = 0; loop_353 < NUM_CELL; loop_353++) begin
         if ({b[1],a[11]}) == loop_353[1:0]) begin
          match_flag_353 = 1'b1;
          addr[353] = loop_353[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_354 = 1'b0;
        addr[354] = 3'b0;
        for (loop_354 = 0; loop_354 < NUM_CELL; loop_354++) begin
         if ({b[2],a[11]}) == loop_354[1:0]) begin
          match_flag_354 = 1'b1;
          addr[354] = loop_354[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_355 = 1'b0;
        addr[355] = 3'b0;
        for (loop_355 = 0; loop_355 < NUM_CELL; loop_355++) begin
         if ({b[3],a[11]}) == loop_355[1:0]) begin
          match_flag_355 = 1'b1;
          addr[355] = loop_355[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_356 = 1'b0;
        addr[356] = 3'b0;
        for (loop_356 = 0; loop_356 < NUM_CELL; loop_356++) begin
         if ({b[4],a[11]}) == loop_356[1:0]) begin
          match_flag_356 = 1'b1;
          addr[356] = loop_356[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_357 = 1'b0;
        addr[357] = 3'b0;
        for (loop_357 = 0; loop_357 < NUM_CELL; loop_357++) begin
         if ({b[5],a[11]}) == loop_357[1:0]) begin
          match_flag_357 = 1'b1;
          addr[357] = loop_357[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_358 = 1'b0;
        addr[358] = 3'b0;
        for (loop_358 = 0; loop_358 < NUM_CELL; loop_358++) begin
         if ({b[6],a[11]}) == loop_358[1:0]) begin
          match_flag_358 = 1'b1;
          addr[358] = loop_358[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_359 = 1'b0;
        addr[359] = 3'b0;
        for (loop_359 = 0; loop_359 < NUM_CELL; loop_359++) begin
         if ({b[7],a[11]}) == loop_359[1:0]) begin
          match_flag_359 = 1'b1;
          addr[359] = loop_359[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_360 = 1'b0;
        addr[360] = 3'b0;
        for (loop_360 = 0; loop_360 < NUM_CELL; loop_360++) begin
         if ({b[8],a[11]}) == loop_360[1:0]) begin
          match_flag_360 = 1'b1;
          addr[360] = loop_360[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_361 = 1'b0;
        addr[361] = 3'b0;
        for (loop_361 = 0; loop_361 < NUM_CELL; loop_361++) begin
         if ({b[9],a[11]}) == loop_361[1:0]) begin
          match_flag_361 = 1'b1;
          addr[361] = loop_361[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_362 = 1'b0;
        addr[362] = 3'b0;
        for (loop_362 = 0; loop_362 < NUM_CELL; loop_362++) begin
         if ({b[10],a[11]}) == loop_362[1:0]) begin
          match_flag_362 = 1'b1;
          addr[362] = loop_362[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_363 = 1'b0;
        addr[363] = 3'b0;
        for (loop_363 = 0; loop_363 < NUM_CELL; loop_363++) begin
         if ({b[11],a[11]}) == loop_363[1:0]) begin
          match_flag_363 = 1'b1;
          addr[363] = loop_363[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_364 = 1'b0;
        addr[364] = 3'b0;
        for (loop_364 = 0; loop_364 < NUM_CELL; loop_364++) begin
         if ({b[12],a[11]}) == loop_364[1:0]) begin
          match_flag_364 = 1'b1;
          addr[364] = loop_364[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_365 = 1'b0;
        addr[365] = 3'b0;
        for (loop_365 = 0; loop_365 < NUM_CELL; loop_365++) begin
         if ({b[13],a[11]}) == loop_365[1:0]) begin
          match_flag_365 = 1'b1;
          addr[365] = loop_365[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_366 = 1'b0;
        addr[366] = 3'b0;
        for (loop_366 = 0; loop_366 < NUM_CELL; loop_366++) begin
         if ({b[14],a[11]}) == loop_366[1:0]) begin
          match_flag_366 = 1'b1;
          addr[366] = loop_366[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_367 = 1'b0;
        addr[367] = 3'b0;
        for (loop_367 = 0; loop_367 < NUM_CELL; loop_367++) begin
         if ({b[15],a[11]}) == loop_367[1:0]) begin
          match_flag_367 = 1'b1;
          addr[367] = loop_367[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_368 = 1'b0;
        addr[368] = 3'b0;
        for (loop_368 = 0; loop_368 < NUM_CELL; loop_368++) begin
         if ({b[16],a[11]}) == loop_368[1:0]) begin
          match_flag_368 = 1'b1;
          addr[368] = loop_368[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_369 = 1'b0;
        addr[369] = 3'b0;
        for (loop_369 = 0; loop_369 < NUM_CELL; loop_369++) begin
         if ({b[17],a[11]}) == loop_369[1:0]) begin
          match_flag_369 = 1'b1;
          addr[369] = loop_369[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_370 = 1'b0;
        addr[370] = 3'b0;
        for (loop_370 = 0; loop_370 < NUM_CELL; loop_370++) begin
         if ({b[18],a[11]}) == loop_370[1:0]) begin
          match_flag_370 = 1'b1;
          addr[370] = loop_370[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_371 = 1'b0;
        addr[371] = 3'b0;
        for (loop_371 = 0; loop_371 < NUM_CELL; loop_371++) begin
         if ({b[19],a[11]}) == loop_371[1:0]) begin
          match_flag_371 = 1'b1;
          addr[371] = loop_371[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_372 = 1'b0;
        addr[372] = 3'b0;
        for (loop_372 = 0; loop_372 < NUM_CELL; loop_372++) begin
         if ({b[20],a[11]}) == loop_372[1:0]) begin
          match_flag_372 = 1'b1;
          addr[372] = loop_372[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_373 = 1'b0;
        addr[373] = 3'b0;
        for (loop_373 = 0; loop_373 < NUM_CELL; loop_373++) begin
         if ({b[21],a[11]}) == loop_373[1:0]) begin
          match_flag_373 = 1'b1;
          addr[373] = loop_373[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_374 = 1'b0;
        addr[374] = 3'b0;
        for (loop_374 = 0; loop_374 < NUM_CELL; loop_374++) begin
         if ({b[22],a[11]}) == loop_374[1:0]) begin
          match_flag_374 = 1'b1;
          addr[374] = loop_374[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_375 = 1'b0;
        addr[375] = 3'b0;
        for (loop_375 = 0; loop_375 < NUM_CELL; loop_375++) begin
         if ({b[23],a[11]}) == loop_375[1:0]) begin
          match_flag_375 = 1'b1;
          addr[375] = loop_375[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_376 = 1'b0;
        addr[376] = 3'b0;
        for (loop_376 = 0; loop_376 < NUM_CELL; loop_376++) begin
         if ({b[24],a[11]}) == loop_376[1:0]) begin
          match_flag_376 = 1'b1;
          addr[376] = loop_376[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_377 = 1'b0;
        addr[377] = 3'b0;
        for (loop_377 = 0; loop_377 < NUM_CELL; loop_377++) begin
         if ({b[25],a[11]}) == loop_377[1:0]) begin
          match_flag_377 = 1'b1;
          addr[377] = loop_377[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_378 = 1'b0;
        addr[378] = 3'b0;
        for (loop_378 = 0; loop_378 < NUM_CELL; loop_378++) begin
         if ({b[26],a[11]}) == loop_378[1:0]) begin
          match_flag_378 = 1'b1;
          addr[378] = loop_378[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_379 = 1'b0;
        addr[379] = 3'b0;
        for (loop_379 = 0; loop_379 < NUM_CELL; loop_379++) begin
         if ({b[27],a[11]}) == loop_379[1:0]) begin
          match_flag_379 = 1'b1;
          addr[379] = loop_379[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_380 = 1'b0;
        addr[380] = 3'b0;
        for (loop_380 = 0; loop_380 < NUM_CELL; loop_380++) begin
         if ({b[28],a[11]}) == loop_380[1:0]) begin
          match_flag_380 = 1'b1;
          addr[380] = loop_380[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_381 = 1'b0;
        addr[381] = 3'b0;
        for (loop_381 = 0; loop_381 < NUM_CELL; loop_381++) begin
         if ({b[29],a[11]}) == loop_381[1:0]) begin
          match_flag_381 = 1'b1;
          addr[381] = loop_381[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_382 = 1'b0;
        addr[382] = 3'b0;
        for (loop_382 = 0; loop_382 < NUM_CELL; loop_382++) begin
         if ({b[30],a[11]}) == loop_382[1:0]) begin
          match_flag_382 = 1'b1;
          addr[382] = loop_382[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_383 = 1'b0;
        addr[383] = 3'b0;
        for (loop_383 = 0; loop_383 < NUM_CELL; loop_383++) begin
         if ({b[31],a[11]}) == loop_383[1:0]) begin
          match_flag_383 = 1'b1;
          addr[383] = loop_383[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_384 = 1'b0;
        addr[384] = 3'b0;
        for (loop_384 = 0; loop_384 < NUM_CELL; loop_384++) begin
         if ({b[0],a[12]}) == loop_384[1:0]) begin
          match_flag_384 = 1'b1;
          addr[384] = loop_384[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_385 = 1'b0;
        addr[385] = 3'b0;
        for (loop_385 = 0; loop_385 < NUM_CELL; loop_385++) begin
         if ({b[1],a[12]}) == loop_385[1:0]) begin
          match_flag_385 = 1'b1;
          addr[385] = loop_385[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_386 = 1'b0;
        addr[386] = 3'b0;
        for (loop_386 = 0; loop_386 < NUM_CELL; loop_386++) begin
         if ({b[2],a[12]}) == loop_386[1:0]) begin
          match_flag_386 = 1'b1;
          addr[386] = loop_386[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_387 = 1'b0;
        addr[387] = 3'b0;
        for (loop_387 = 0; loop_387 < NUM_CELL; loop_387++) begin
         if ({b[3],a[12]}) == loop_387[1:0]) begin
          match_flag_387 = 1'b1;
          addr[387] = loop_387[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_388 = 1'b0;
        addr[388] = 3'b0;
        for (loop_388 = 0; loop_388 < NUM_CELL; loop_388++) begin
         if ({b[4],a[12]}) == loop_388[1:0]) begin
          match_flag_388 = 1'b1;
          addr[388] = loop_388[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_389 = 1'b0;
        addr[389] = 3'b0;
        for (loop_389 = 0; loop_389 < NUM_CELL; loop_389++) begin
         if ({b[5],a[12]}) == loop_389[1:0]) begin
          match_flag_389 = 1'b1;
          addr[389] = loop_389[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_390 = 1'b0;
        addr[390] = 3'b0;
        for (loop_390 = 0; loop_390 < NUM_CELL; loop_390++) begin
         if ({b[6],a[12]}) == loop_390[1:0]) begin
          match_flag_390 = 1'b1;
          addr[390] = loop_390[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_391 = 1'b0;
        addr[391] = 3'b0;
        for (loop_391 = 0; loop_391 < NUM_CELL; loop_391++) begin
         if ({b[7],a[12]}) == loop_391[1:0]) begin
          match_flag_391 = 1'b1;
          addr[391] = loop_391[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_392 = 1'b0;
        addr[392] = 3'b0;
        for (loop_392 = 0; loop_392 < NUM_CELL; loop_392++) begin
         if ({b[8],a[12]}) == loop_392[1:0]) begin
          match_flag_392 = 1'b1;
          addr[392] = loop_392[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_393 = 1'b0;
        addr[393] = 3'b0;
        for (loop_393 = 0; loop_393 < NUM_CELL; loop_393++) begin
         if ({b[9],a[12]}) == loop_393[1:0]) begin
          match_flag_393 = 1'b1;
          addr[393] = loop_393[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_394 = 1'b0;
        addr[394] = 3'b0;
        for (loop_394 = 0; loop_394 < NUM_CELL; loop_394++) begin
         if ({b[10],a[12]}) == loop_394[1:0]) begin
          match_flag_394 = 1'b1;
          addr[394] = loop_394[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_395 = 1'b0;
        addr[395] = 3'b0;
        for (loop_395 = 0; loop_395 < NUM_CELL; loop_395++) begin
         if ({b[11],a[12]}) == loop_395[1:0]) begin
          match_flag_395 = 1'b1;
          addr[395] = loop_395[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_396 = 1'b0;
        addr[396] = 3'b0;
        for (loop_396 = 0; loop_396 < NUM_CELL; loop_396++) begin
         if ({b[12],a[12]}) == loop_396[1:0]) begin
          match_flag_396 = 1'b1;
          addr[396] = loop_396[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_397 = 1'b0;
        addr[397] = 3'b0;
        for (loop_397 = 0; loop_397 < NUM_CELL; loop_397++) begin
         if ({b[13],a[12]}) == loop_397[1:0]) begin
          match_flag_397 = 1'b1;
          addr[397] = loop_397[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_398 = 1'b0;
        addr[398] = 3'b0;
        for (loop_398 = 0; loop_398 < NUM_CELL; loop_398++) begin
         if ({b[14],a[12]}) == loop_398[1:0]) begin
          match_flag_398 = 1'b1;
          addr[398] = loop_398[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_399 = 1'b0;
        addr[399] = 3'b0;
        for (loop_399 = 0; loop_399 < NUM_CELL; loop_399++) begin
         if ({b[15],a[12]}) == loop_399[1:0]) begin
          match_flag_399 = 1'b1;
          addr[399] = loop_399[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_400 = 1'b0;
        addr[400] = 3'b0;
        for (loop_400 = 0; loop_400 < NUM_CELL; loop_400++) begin
         if ({b[16],a[12]}) == loop_400[1:0]) begin
          match_flag_400 = 1'b1;
          addr[400] = loop_400[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_401 = 1'b0;
        addr[401] = 3'b0;
        for (loop_401 = 0; loop_401 < NUM_CELL; loop_401++) begin
         if ({b[17],a[12]}) == loop_401[1:0]) begin
          match_flag_401 = 1'b1;
          addr[401] = loop_401[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_402 = 1'b0;
        addr[402] = 3'b0;
        for (loop_402 = 0; loop_402 < NUM_CELL; loop_402++) begin
         if ({b[18],a[12]}) == loop_402[1:0]) begin
          match_flag_402 = 1'b1;
          addr[402] = loop_402[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_403 = 1'b0;
        addr[403] = 3'b0;
        for (loop_403 = 0; loop_403 < NUM_CELL; loop_403++) begin
         if ({b[19],a[12]}) == loop_403[1:0]) begin
          match_flag_403 = 1'b1;
          addr[403] = loop_403[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_404 = 1'b0;
        addr[404] = 3'b0;
        for (loop_404 = 0; loop_404 < NUM_CELL; loop_404++) begin
         if ({b[20],a[12]}) == loop_404[1:0]) begin
          match_flag_404 = 1'b1;
          addr[404] = loop_404[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_405 = 1'b0;
        addr[405] = 3'b0;
        for (loop_405 = 0; loop_405 < NUM_CELL; loop_405++) begin
         if ({b[21],a[12]}) == loop_405[1:0]) begin
          match_flag_405 = 1'b1;
          addr[405] = loop_405[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_406 = 1'b0;
        addr[406] = 3'b0;
        for (loop_406 = 0; loop_406 < NUM_CELL; loop_406++) begin
         if ({b[22],a[12]}) == loop_406[1:0]) begin
          match_flag_406 = 1'b1;
          addr[406] = loop_406[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_407 = 1'b0;
        addr[407] = 3'b0;
        for (loop_407 = 0; loop_407 < NUM_CELL; loop_407++) begin
         if ({b[23],a[12]}) == loop_407[1:0]) begin
          match_flag_407 = 1'b1;
          addr[407] = loop_407[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_408 = 1'b0;
        addr[408] = 3'b0;
        for (loop_408 = 0; loop_408 < NUM_CELL; loop_408++) begin
         if ({b[24],a[12]}) == loop_408[1:0]) begin
          match_flag_408 = 1'b1;
          addr[408] = loop_408[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_409 = 1'b0;
        addr[409] = 3'b0;
        for (loop_409 = 0; loop_409 < NUM_CELL; loop_409++) begin
         if ({b[25],a[12]}) == loop_409[1:0]) begin
          match_flag_409 = 1'b1;
          addr[409] = loop_409[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_410 = 1'b0;
        addr[410] = 3'b0;
        for (loop_410 = 0; loop_410 < NUM_CELL; loop_410++) begin
         if ({b[26],a[12]}) == loop_410[1:0]) begin
          match_flag_410 = 1'b1;
          addr[410] = loop_410[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_411 = 1'b0;
        addr[411] = 3'b0;
        for (loop_411 = 0; loop_411 < NUM_CELL; loop_411++) begin
         if ({b[27],a[12]}) == loop_411[1:0]) begin
          match_flag_411 = 1'b1;
          addr[411] = loop_411[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_412 = 1'b0;
        addr[412] = 3'b0;
        for (loop_412 = 0; loop_412 < NUM_CELL; loop_412++) begin
         if ({b[28],a[12]}) == loop_412[1:0]) begin
          match_flag_412 = 1'b1;
          addr[412] = loop_412[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_413 = 1'b0;
        addr[413] = 3'b0;
        for (loop_413 = 0; loop_413 < NUM_CELL; loop_413++) begin
         if ({b[29],a[12]}) == loop_413[1:0]) begin
          match_flag_413 = 1'b1;
          addr[413] = loop_413[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_414 = 1'b0;
        addr[414] = 3'b0;
        for (loop_414 = 0; loop_414 < NUM_CELL; loop_414++) begin
         if ({b[30],a[12]}) == loop_414[1:0]) begin
          match_flag_414 = 1'b1;
          addr[414] = loop_414[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_415 = 1'b0;
        addr[415] = 3'b0;
        for (loop_415 = 0; loop_415 < NUM_CELL; loop_415++) begin
         if ({b[31],a[12]}) == loop_415[1:0]) begin
          match_flag_415 = 1'b1;
          addr[415] = loop_415[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_416 = 1'b0;
        addr[416] = 3'b0;
        for (loop_416 = 0; loop_416 < NUM_CELL; loop_416++) begin
         if ({b[0],a[13]}) == loop_416[1:0]) begin
          match_flag_416 = 1'b1;
          addr[416] = loop_416[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_417 = 1'b0;
        addr[417] = 3'b0;
        for (loop_417 = 0; loop_417 < NUM_CELL; loop_417++) begin
         if ({b[1],a[13]}) == loop_417[1:0]) begin
          match_flag_417 = 1'b1;
          addr[417] = loop_417[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_418 = 1'b0;
        addr[418] = 3'b0;
        for (loop_418 = 0; loop_418 < NUM_CELL; loop_418++) begin
         if ({b[2],a[13]}) == loop_418[1:0]) begin
          match_flag_418 = 1'b1;
          addr[418] = loop_418[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_419 = 1'b0;
        addr[419] = 3'b0;
        for (loop_419 = 0; loop_419 < NUM_CELL; loop_419++) begin
         if ({b[3],a[13]}) == loop_419[1:0]) begin
          match_flag_419 = 1'b1;
          addr[419] = loop_419[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_420 = 1'b0;
        addr[420] = 3'b0;
        for (loop_420 = 0; loop_420 < NUM_CELL; loop_420++) begin
         if ({b[4],a[13]}) == loop_420[1:0]) begin
          match_flag_420 = 1'b1;
          addr[420] = loop_420[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_421 = 1'b0;
        addr[421] = 3'b0;
        for (loop_421 = 0; loop_421 < NUM_CELL; loop_421++) begin
         if ({b[5],a[13]}) == loop_421[1:0]) begin
          match_flag_421 = 1'b1;
          addr[421] = loop_421[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_422 = 1'b0;
        addr[422] = 3'b0;
        for (loop_422 = 0; loop_422 < NUM_CELL; loop_422++) begin
         if ({b[6],a[13]}) == loop_422[1:0]) begin
          match_flag_422 = 1'b1;
          addr[422] = loop_422[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_423 = 1'b0;
        addr[423] = 3'b0;
        for (loop_423 = 0; loop_423 < NUM_CELL; loop_423++) begin
         if ({b[7],a[13]}) == loop_423[1:0]) begin
          match_flag_423 = 1'b1;
          addr[423] = loop_423[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_424 = 1'b0;
        addr[424] = 3'b0;
        for (loop_424 = 0; loop_424 < NUM_CELL; loop_424++) begin
         if ({b[8],a[13]}) == loop_424[1:0]) begin
          match_flag_424 = 1'b1;
          addr[424] = loop_424[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_425 = 1'b0;
        addr[425] = 3'b0;
        for (loop_425 = 0; loop_425 < NUM_CELL; loop_425++) begin
         if ({b[9],a[13]}) == loop_425[1:0]) begin
          match_flag_425 = 1'b1;
          addr[425] = loop_425[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_426 = 1'b0;
        addr[426] = 3'b0;
        for (loop_426 = 0; loop_426 < NUM_CELL; loop_426++) begin
         if ({b[10],a[13]}) == loop_426[1:0]) begin
          match_flag_426 = 1'b1;
          addr[426] = loop_426[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_427 = 1'b0;
        addr[427] = 3'b0;
        for (loop_427 = 0; loop_427 < NUM_CELL; loop_427++) begin
         if ({b[11],a[13]}) == loop_427[1:0]) begin
          match_flag_427 = 1'b1;
          addr[427] = loop_427[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_428 = 1'b0;
        addr[428] = 3'b0;
        for (loop_428 = 0; loop_428 < NUM_CELL; loop_428++) begin
         if ({b[12],a[13]}) == loop_428[1:0]) begin
          match_flag_428 = 1'b1;
          addr[428] = loop_428[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_429 = 1'b0;
        addr[429] = 3'b0;
        for (loop_429 = 0; loop_429 < NUM_CELL; loop_429++) begin
         if ({b[13],a[13]}) == loop_429[1:0]) begin
          match_flag_429 = 1'b1;
          addr[429] = loop_429[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_430 = 1'b0;
        addr[430] = 3'b0;
        for (loop_430 = 0; loop_430 < NUM_CELL; loop_430++) begin
         if ({b[14],a[13]}) == loop_430[1:0]) begin
          match_flag_430 = 1'b1;
          addr[430] = loop_430[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_431 = 1'b0;
        addr[431] = 3'b0;
        for (loop_431 = 0; loop_431 < NUM_CELL; loop_431++) begin
         if ({b[15],a[13]}) == loop_431[1:0]) begin
          match_flag_431 = 1'b1;
          addr[431] = loop_431[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_432 = 1'b0;
        addr[432] = 3'b0;
        for (loop_432 = 0; loop_432 < NUM_CELL; loop_432++) begin
         if ({b[16],a[13]}) == loop_432[1:0]) begin
          match_flag_432 = 1'b1;
          addr[432] = loop_432[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_433 = 1'b0;
        addr[433] = 3'b0;
        for (loop_433 = 0; loop_433 < NUM_CELL; loop_433++) begin
         if ({b[17],a[13]}) == loop_433[1:0]) begin
          match_flag_433 = 1'b1;
          addr[433] = loop_433[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_434 = 1'b0;
        addr[434] = 3'b0;
        for (loop_434 = 0; loop_434 < NUM_CELL; loop_434++) begin
         if ({b[18],a[13]}) == loop_434[1:0]) begin
          match_flag_434 = 1'b1;
          addr[434] = loop_434[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_435 = 1'b0;
        addr[435] = 3'b0;
        for (loop_435 = 0; loop_435 < NUM_CELL; loop_435++) begin
         if ({b[19],a[13]}) == loop_435[1:0]) begin
          match_flag_435 = 1'b1;
          addr[435] = loop_435[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_436 = 1'b0;
        addr[436] = 3'b0;
        for (loop_436 = 0; loop_436 < NUM_CELL; loop_436++) begin
         if ({b[20],a[13]}) == loop_436[1:0]) begin
          match_flag_436 = 1'b1;
          addr[436] = loop_436[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_437 = 1'b0;
        addr[437] = 3'b0;
        for (loop_437 = 0; loop_437 < NUM_CELL; loop_437++) begin
         if ({b[21],a[13]}) == loop_437[1:0]) begin
          match_flag_437 = 1'b1;
          addr[437] = loop_437[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_438 = 1'b0;
        addr[438] = 3'b0;
        for (loop_438 = 0; loop_438 < NUM_CELL; loop_438++) begin
         if ({b[22],a[13]}) == loop_438[1:0]) begin
          match_flag_438 = 1'b1;
          addr[438] = loop_438[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_439 = 1'b0;
        addr[439] = 3'b0;
        for (loop_439 = 0; loop_439 < NUM_CELL; loop_439++) begin
         if ({b[23],a[13]}) == loop_439[1:0]) begin
          match_flag_439 = 1'b1;
          addr[439] = loop_439[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_440 = 1'b0;
        addr[440] = 3'b0;
        for (loop_440 = 0; loop_440 < NUM_CELL; loop_440++) begin
         if ({b[24],a[13]}) == loop_440[1:0]) begin
          match_flag_440 = 1'b1;
          addr[440] = loop_440[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_441 = 1'b0;
        addr[441] = 3'b0;
        for (loop_441 = 0; loop_441 < NUM_CELL; loop_441++) begin
         if ({b[25],a[13]}) == loop_441[1:0]) begin
          match_flag_441 = 1'b1;
          addr[441] = loop_441[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_442 = 1'b0;
        addr[442] = 3'b0;
        for (loop_442 = 0; loop_442 < NUM_CELL; loop_442++) begin
         if ({b[26],a[13]}) == loop_442[1:0]) begin
          match_flag_442 = 1'b1;
          addr[442] = loop_442[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_443 = 1'b0;
        addr[443] = 3'b0;
        for (loop_443 = 0; loop_443 < NUM_CELL; loop_443++) begin
         if ({b[27],a[13]}) == loop_443[1:0]) begin
          match_flag_443 = 1'b1;
          addr[443] = loop_443[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_444 = 1'b0;
        addr[444] = 3'b0;
        for (loop_444 = 0; loop_444 < NUM_CELL; loop_444++) begin
         if ({b[28],a[13]}) == loop_444[1:0]) begin
          match_flag_444 = 1'b1;
          addr[444] = loop_444[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_445 = 1'b0;
        addr[445] = 3'b0;
        for (loop_445 = 0; loop_445 < NUM_CELL; loop_445++) begin
         if ({b[29],a[13]}) == loop_445[1:0]) begin
          match_flag_445 = 1'b1;
          addr[445] = loop_445[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_446 = 1'b0;
        addr[446] = 3'b0;
        for (loop_446 = 0; loop_446 < NUM_CELL; loop_446++) begin
         if ({b[30],a[13]}) == loop_446[1:0]) begin
          match_flag_446 = 1'b1;
          addr[446] = loop_446[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_447 = 1'b0;
        addr[447] = 3'b0;
        for (loop_447 = 0; loop_447 < NUM_CELL; loop_447++) begin
         if ({b[31],a[13]}) == loop_447[1:0]) begin
          match_flag_447 = 1'b1;
          addr[447] = loop_447[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_448 = 1'b0;
        addr[448] = 3'b0;
        for (loop_448 = 0; loop_448 < NUM_CELL; loop_448++) begin
         if ({b[0],a[14]}) == loop_448[1:0]) begin
          match_flag_448 = 1'b1;
          addr[448] = loop_448[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_449 = 1'b0;
        addr[449] = 3'b0;
        for (loop_449 = 0; loop_449 < NUM_CELL; loop_449++) begin
         if ({b[1],a[14]}) == loop_449[1:0]) begin
          match_flag_449 = 1'b1;
          addr[449] = loop_449[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_450 = 1'b0;
        addr[450] = 3'b0;
        for (loop_450 = 0; loop_450 < NUM_CELL; loop_450++) begin
         if ({b[2],a[14]}) == loop_450[1:0]) begin
          match_flag_450 = 1'b1;
          addr[450] = loop_450[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_451 = 1'b0;
        addr[451] = 3'b0;
        for (loop_451 = 0; loop_451 < NUM_CELL; loop_451++) begin
         if ({b[3],a[14]}) == loop_451[1:0]) begin
          match_flag_451 = 1'b1;
          addr[451] = loop_451[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_452 = 1'b0;
        addr[452] = 3'b0;
        for (loop_452 = 0; loop_452 < NUM_CELL; loop_452++) begin
         if ({b[4],a[14]}) == loop_452[1:0]) begin
          match_flag_452 = 1'b1;
          addr[452] = loop_452[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_453 = 1'b0;
        addr[453] = 3'b0;
        for (loop_453 = 0; loop_453 < NUM_CELL; loop_453++) begin
         if ({b[5],a[14]}) == loop_453[1:0]) begin
          match_flag_453 = 1'b1;
          addr[453] = loop_453[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_454 = 1'b0;
        addr[454] = 3'b0;
        for (loop_454 = 0; loop_454 < NUM_CELL; loop_454++) begin
         if ({b[6],a[14]}) == loop_454[1:0]) begin
          match_flag_454 = 1'b1;
          addr[454] = loop_454[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_455 = 1'b0;
        addr[455] = 3'b0;
        for (loop_455 = 0; loop_455 < NUM_CELL; loop_455++) begin
         if ({b[7],a[14]}) == loop_455[1:0]) begin
          match_flag_455 = 1'b1;
          addr[455] = loop_455[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_456 = 1'b0;
        addr[456] = 3'b0;
        for (loop_456 = 0; loop_456 < NUM_CELL; loop_456++) begin
         if ({b[8],a[14]}) == loop_456[1:0]) begin
          match_flag_456 = 1'b1;
          addr[456] = loop_456[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_457 = 1'b0;
        addr[457] = 3'b0;
        for (loop_457 = 0; loop_457 < NUM_CELL; loop_457++) begin
         if ({b[9],a[14]}) == loop_457[1:0]) begin
          match_flag_457 = 1'b1;
          addr[457] = loop_457[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_458 = 1'b0;
        addr[458] = 3'b0;
        for (loop_458 = 0; loop_458 < NUM_CELL; loop_458++) begin
         if ({b[10],a[14]}) == loop_458[1:0]) begin
          match_flag_458 = 1'b1;
          addr[458] = loop_458[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_459 = 1'b0;
        addr[459] = 3'b0;
        for (loop_459 = 0; loop_459 < NUM_CELL; loop_459++) begin
         if ({b[11],a[14]}) == loop_459[1:0]) begin
          match_flag_459 = 1'b1;
          addr[459] = loop_459[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_460 = 1'b0;
        addr[460] = 3'b0;
        for (loop_460 = 0; loop_460 < NUM_CELL; loop_460++) begin
         if ({b[12],a[14]}) == loop_460[1:0]) begin
          match_flag_460 = 1'b1;
          addr[460] = loop_460[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_461 = 1'b0;
        addr[461] = 3'b0;
        for (loop_461 = 0; loop_461 < NUM_CELL; loop_461++) begin
         if ({b[13],a[14]}) == loop_461[1:0]) begin
          match_flag_461 = 1'b1;
          addr[461] = loop_461[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_462 = 1'b0;
        addr[462] = 3'b0;
        for (loop_462 = 0; loop_462 < NUM_CELL; loop_462++) begin
         if ({b[14],a[14]}) == loop_462[1:0]) begin
          match_flag_462 = 1'b1;
          addr[462] = loop_462[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_463 = 1'b0;
        addr[463] = 3'b0;
        for (loop_463 = 0; loop_463 < NUM_CELL; loop_463++) begin
         if ({b[15],a[14]}) == loop_463[1:0]) begin
          match_flag_463 = 1'b1;
          addr[463] = loop_463[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_464 = 1'b0;
        addr[464] = 3'b0;
        for (loop_464 = 0; loop_464 < NUM_CELL; loop_464++) begin
         if ({b[16],a[14]}) == loop_464[1:0]) begin
          match_flag_464 = 1'b1;
          addr[464] = loop_464[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_465 = 1'b0;
        addr[465] = 3'b0;
        for (loop_465 = 0; loop_465 < NUM_CELL; loop_465++) begin
         if ({b[17],a[14]}) == loop_465[1:0]) begin
          match_flag_465 = 1'b1;
          addr[465] = loop_465[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_466 = 1'b0;
        addr[466] = 3'b0;
        for (loop_466 = 0; loop_466 < NUM_CELL; loop_466++) begin
         if ({b[18],a[14]}) == loop_466[1:0]) begin
          match_flag_466 = 1'b1;
          addr[466] = loop_466[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_467 = 1'b0;
        addr[467] = 3'b0;
        for (loop_467 = 0; loop_467 < NUM_CELL; loop_467++) begin
         if ({b[19],a[14]}) == loop_467[1:0]) begin
          match_flag_467 = 1'b1;
          addr[467] = loop_467[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_468 = 1'b0;
        addr[468] = 3'b0;
        for (loop_468 = 0; loop_468 < NUM_CELL; loop_468++) begin
         if ({b[20],a[14]}) == loop_468[1:0]) begin
          match_flag_468 = 1'b1;
          addr[468] = loop_468[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_469 = 1'b0;
        addr[469] = 3'b0;
        for (loop_469 = 0; loop_469 < NUM_CELL; loop_469++) begin
         if ({b[21],a[14]}) == loop_469[1:0]) begin
          match_flag_469 = 1'b1;
          addr[469] = loop_469[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_470 = 1'b0;
        addr[470] = 3'b0;
        for (loop_470 = 0; loop_470 < NUM_CELL; loop_470++) begin
         if ({b[22],a[14]}) == loop_470[1:0]) begin
          match_flag_470 = 1'b1;
          addr[470] = loop_470[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_471 = 1'b0;
        addr[471] = 3'b0;
        for (loop_471 = 0; loop_471 < NUM_CELL; loop_471++) begin
         if ({b[23],a[14]}) == loop_471[1:0]) begin
          match_flag_471 = 1'b1;
          addr[471] = loop_471[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_472 = 1'b0;
        addr[472] = 3'b0;
        for (loop_472 = 0; loop_472 < NUM_CELL; loop_472++) begin
         if ({b[24],a[14]}) == loop_472[1:0]) begin
          match_flag_472 = 1'b1;
          addr[472] = loop_472[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_473 = 1'b0;
        addr[473] = 3'b0;
        for (loop_473 = 0; loop_473 < NUM_CELL; loop_473++) begin
         if ({b[25],a[14]}) == loop_473[1:0]) begin
          match_flag_473 = 1'b1;
          addr[473] = loop_473[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_474 = 1'b0;
        addr[474] = 3'b0;
        for (loop_474 = 0; loop_474 < NUM_CELL; loop_474++) begin
         if ({b[26],a[14]}) == loop_474[1:0]) begin
          match_flag_474 = 1'b1;
          addr[474] = loop_474[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_475 = 1'b0;
        addr[475] = 3'b0;
        for (loop_475 = 0; loop_475 < NUM_CELL; loop_475++) begin
         if ({b[27],a[14]}) == loop_475[1:0]) begin
          match_flag_475 = 1'b1;
          addr[475] = loop_475[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_476 = 1'b0;
        addr[476] = 3'b0;
        for (loop_476 = 0; loop_476 < NUM_CELL; loop_476++) begin
         if ({b[28],a[14]}) == loop_476[1:0]) begin
          match_flag_476 = 1'b1;
          addr[476] = loop_476[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_477 = 1'b0;
        addr[477] = 3'b0;
        for (loop_477 = 0; loop_477 < NUM_CELL; loop_477++) begin
         if ({b[29],a[14]}) == loop_477[1:0]) begin
          match_flag_477 = 1'b1;
          addr[477] = loop_477[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_478 = 1'b0;
        addr[478] = 3'b0;
        for (loop_478 = 0; loop_478 < NUM_CELL; loop_478++) begin
         if ({b[30],a[14]}) == loop_478[1:0]) begin
          match_flag_478 = 1'b1;
          addr[478] = loop_478[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_479 = 1'b0;
        addr[479] = 3'b0;
        for (loop_479 = 0; loop_479 < NUM_CELL; loop_479++) begin
         if ({b[31],a[14]}) == loop_479[1:0]) begin
          match_flag_479 = 1'b1;
          addr[479] = loop_479[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_480 = 1'b0;
        addr[480] = 3'b0;
        for (loop_480 = 0; loop_480 < NUM_CELL; loop_480++) begin
         if ({b[0],a[15]}) == loop_480[1:0]) begin
          match_flag_480 = 1'b1;
          addr[480] = loop_480[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_481 = 1'b0;
        addr[481] = 3'b0;
        for (loop_481 = 0; loop_481 < NUM_CELL; loop_481++) begin
         if ({b[1],a[15]}) == loop_481[1:0]) begin
          match_flag_481 = 1'b1;
          addr[481] = loop_481[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_482 = 1'b0;
        addr[482] = 3'b0;
        for (loop_482 = 0; loop_482 < NUM_CELL; loop_482++) begin
         if ({b[2],a[15]}) == loop_482[1:0]) begin
          match_flag_482 = 1'b1;
          addr[482] = loop_482[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_483 = 1'b0;
        addr[483] = 3'b0;
        for (loop_483 = 0; loop_483 < NUM_CELL; loop_483++) begin
         if ({b[3],a[15]}) == loop_483[1:0]) begin
          match_flag_483 = 1'b1;
          addr[483] = loop_483[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_484 = 1'b0;
        addr[484] = 3'b0;
        for (loop_484 = 0; loop_484 < NUM_CELL; loop_484++) begin
         if ({b[4],a[15]}) == loop_484[1:0]) begin
          match_flag_484 = 1'b1;
          addr[484] = loop_484[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_485 = 1'b0;
        addr[485] = 3'b0;
        for (loop_485 = 0; loop_485 < NUM_CELL; loop_485++) begin
         if ({b[5],a[15]}) == loop_485[1:0]) begin
          match_flag_485 = 1'b1;
          addr[485] = loop_485[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_486 = 1'b0;
        addr[486] = 3'b0;
        for (loop_486 = 0; loop_486 < NUM_CELL; loop_486++) begin
         if ({b[6],a[15]}) == loop_486[1:0]) begin
          match_flag_486 = 1'b1;
          addr[486] = loop_486[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_487 = 1'b0;
        addr[487] = 3'b0;
        for (loop_487 = 0; loop_487 < NUM_CELL; loop_487++) begin
         if ({b[7],a[15]}) == loop_487[1:0]) begin
          match_flag_487 = 1'b1;
          addr[487] = loop_487[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_488 = 1'b0;
        addr[488] = 3'b0;
        for (loop_488 = 0; loop_488 < NUM_CELL; loop_488++) begin
         if ({b[8],a[15]}) == loop_488[1:0]) begin
          match_flag_488 = 1'b1;
          addr[488] = loop_488[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_489 = 1'b0;
        addr[489] = 3'b0;
        for (loop_489 = 0; loop_489 < NUM_CELL; loop_489++) begin
         if ({b[9],a[15]}) == loop_489[1:0]) begin
          match_flag_489 = 1'b1;
          addr[489] = loop_489[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_490 = 1'b0;
        addr[490] = 3'b0;
        for (loop_490 = 0; loop_490 < NUM_CELL; loop_490++) begin
         if ({b[10],a[15]}) == loop_490[1:0]) begin
          match_flag_490 = 1'b1;
          addr[490] = loop_490[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_491 = 1'b0;
        addr[491] = 3'b0;
        for (loop_491 = 0; loop_491 < NUM_CELL; loop_491++) begin
         if ({b[11],a[15]}) == loop_491[1:0]) begin
          match_flag_491 = 1'b1;
          addr[491] = loop_491[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_492 = 1'b0;
        addr[492] = 3'b0;
        for (loop_492 = 0; loop_492 < NUM_CELL; loop_492++) begin
         if ({b[12],a[15]}) == loop_492[1:0]) begin
          match_flag_492 = 1'b1;
          addr[492] = loop_492[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_493 = 1'b0;
        addr[493] = 3'b0;
        for (loop_493 = 0; loop_493 < NUM_CELL; loop_493++) begin
         if ({b[13],a[15]}) == loop_493[1:0]) begin
          match_flag_493 = 1'b1;
          addr[493] = loop_493[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_494 = 1'b0;
        addr[494] = 3'b0;
        for (loop_494 = 0; loop_494 < NUM_CELL; loop_494++) begin
         if ({b[14],a[15]}) == loop_494[1:0]) begin
          match_flag_494 = 1'b1;
          addr[494] = loop_494[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_495 = 1'b0;
        addr[495] = 3'b0;
        for (loop_495 = 0; loop_495 < NUM_CELL; loop_495++) begin
         if ({b[15],a[15]}) == loop_495[1:0]) begin
          match_flag_495 = 1'b1;
          addr[495] = loop_495[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_496 = 1'b0;
        addr[496] = 3'b0;
        for (loop_496 = 0; loop_496 < NUM_CELL; loop_496++) begin
         if ({b[16],a[15]}) == loop_496[1:0]) begin
          match_flag_496 = 1'b1;
          addr[496] = loop_496[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_497 = 1'b0;
        addr[497] = 3'b0;
        for (loop_497 = 0; loop_497 < NUM_CELL; loop_497++) begin
         if ({b[17],a[15]}) == loop_497[1:0]) begin
          match_flag_497 = 1'b1;
          addr[497] = loop_497[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_498 = 1'b0;
        addr[498] = 3'b0;
        for (loop_498 = 0; loop_498 < NUM_CELL; loop_498++) begin
         if ({b[18],a[15]}) == loop_498[1:0]) begin
          match_flag_498 = 1'b1;
          addr[498] = loop_498[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_499 = 1'b0;
        addr[499] = 3'b0;
        for (loop_499 = 0; loop_499 < NUM_CELL; loop_499++) begin
         if ({b[19],a[15]}) == loop_499[1:0]) begin
          match_flag_499 = 1'b1;
          addr[499] = loop_499[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_500 = 1'b0;
        addr[500] = 3'b0;
        for (loop_500 = 0; loop_500 < NUM_CELL; loop_500++) begin
         if ({b[20],a[15]}) == loop_500[1:0]) begin
          match_flag_500 = 1'b1;
          addr[500] = loop_500[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_501 = 1'b0;
        addr[501] = 3'b0;
        for (loop_501 = 0; loop_501 < NUM_CELL; loop_501++) begin
         if ({b[21],a[15]}) == loop_501[1:0]) begin
          match_flag_501 = 1'b1;
          addr[501] = loop_501[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_502 = 1'b0;
        addr[502] = 3'b0;
        for (loop_502 = 0; loop_502 < NUM_CELL; loop_502++) begin
         if ({b[22],a[15]}) == loop_502[1:0]) begin
          match_flag_502 = 1'b1;
          addr[502] = loop_502[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_503 = 1'b0;
        addr[503] = 3'b0;
        for (loop_503 = 0; loop_503 < NUM_CELL; loop_503++) begin
         if ({b[23],a[15]}) == loop_503[1:0]) begin
          match_flag_503 = 1'b1;
          addr[503] = loop_503[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_504 = 1'b0;
        addr[504] = 3'b0;
        for (loop_504 = 0; loop_504 < NUM_CELL; loop_504++) begin
         if ({b[24],a[15]}) == loop_504[1:0]) begin
          match_flag_504 = 1'b1;
          addr[504] = loop_504[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_505 = 1'b0;
        addr[505] = 3'b0;
        for (loop_505 = 0; loop_505 < NUM_CELL; loop_505++) begin
         if ({b[25],a[15]}) == loop_505[1:0]) begin
          match_flag_505 = 1'b1;
          addr[505] = loop_505[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_506 = 1'b0;
        addr[506] = 3'b0;
        for (loop_506 = 0; loop_506 < NUM_CELL; loop_506++) begin
         if ({b[26],a[15]}) == loop_506[1:0]) begin
          match_flag_506 = 1'b1;
          addr[506] = loop_506[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_507 = 1'b0;
        addr[507] = 3'b0;
        for (loop_507 = 0; loop_507 < NUM_CELL; loop_507++) begin
         if ({b[27],a[15]}) == loop_507[1:0]) begin
          match_flag_507 = 1'b1;
          addr[507] = loop_507[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_508 = 1'b0;
        addr[508] = 3'b0;
        for (loop_508 = 0; loop_508 < NUM_CELL; loop_508++) begin
         if ({b[28],a[15]}) == loop_508[1:0]) begin
          match_flag_508 = 1'b1;
          addr[508] = loop_508[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_509 = 1'b0;
        addr[509] = 3'b0;
        for (loop_509 = 0; loop_509 < NUM_CELL; loop_509++) begin
         if ({b[29],a[15]}) == loop_509[1:0]) begin
          match_flag_509 = 1'b1;
          addr[509] = loop_509[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_510 = 1'b0;
        addr[510] = 3'b0;
        for (loop_510 = 0; loop_510 < NUM_CELL; loop_510++) begin
         if ({b[30],a[15]}) == loop_510[1:0]) begin
          match_flag_510 = 1'b1;
          addr[510] = loop_510[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_511 = 1'b0;
        addr[511] = 3'b0;
        for (loop_511 = 0; loop_511 < NUM_CELL; loop_511++) begin
         if ({b[31],a[15]}) == loop_511[1:0]) begin
          match_flag_511 = 1'b1;
          addr[511] = loop_511[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_512 = 1'b0;
        addr[512] = 3'b0;
        for (loop_512 = 0; loop_512 < NUM_CELL; loop_512++) begin
         if ({b[0],a[16]}) == loop_512[1:0]) begin
          match_flag_512 = 1'b1;
          addr[512] = loop_512[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_513 = 1'b0;
        addr[513] = 3'b0;
        for (loop_513 = 0; loop_513 < NUM_CELL; loop_513++) begin
         if ({b[1],a[16]}) == loop_513[1:0]) begin
          match_flag_513 = 1'b1;
          addr[513] = loop_513[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_514 = 1'b0;
        addr[514] = 3'b0;
        for (loop_514 = 0; loop_514 < NUM_CELL; loop_514++) begin
         if ({b[2],a[16]}) == loop_514[1:0]) begin
          match_flag_514 = 1'b1;
          addr[514] = loop_514[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_515 = 1'b0;
        addr[515] = 3'b0;
        for (loop_515 = 0; loop_515 < NUM_CELL; loop_515++) begin
         if ({b[3],a[16]}) == loop_515[1:0]) begin
          match_flag_515 = 1'b1;
          addr[515] = loop_515[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_516 = 1'b0;
        addr[516] = 3'b0;
        for (loop_516 = 0; loop_516 < NUM_CELL; loop_516++) begin
         if ({b[4],a[16]}) == loop_516[1:0]) begin
          match_flag_516 = 1'b1;
          addr[516] = loop_516[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_517 = 1'b0;
        addr[517] = 3'b0;
        for (loop_517 = 0; loop_517 < NUM_CELL; loop_517++) begin
         if ({b[5],a[16]}) == loop_517[1:0]) begin
          match_flag_517 = 1'b1;
          addr[517] = loop_517[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_518 = 1'b0;
        addr[518] = 3'b0;
        for (loop_518 = 0; loop_518 < NUM_CELL; loop_518++) begin
         if ({b[6],a[16]}) == loop_518[1:0]) begin
          match_flag_518 = 1'b1;
          addr[518] = loop_518[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_519 = 1'b0;
        addr[519] = 3'b0;
        for (loop_519 = 0; loop_519 < NUM_CELL; loop_519++) begin
         if ({b[7],a[16]}) == loop_519[1:0]) begin
          match_flag_519 = 1'b1;
          addr[519] = loop_519[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_520 = 1'b0;
        addr[520] = 3'b0;
        for (loop_520 = 0; loop_520 < NUM_CELL; loop_520++) begin
         if ({b[8],a[16]}) == loop_520[1:0]) begin
          match_flag_520 = 1'b1;
          addr[520] = loop_520[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_521 = 1'b0;
        addr[521] = 3'b0;
        for (loop_521 = 0; loop_521 < NUM_CELL; loop_521++) begin
         if ({b[9],a[16]}) == loop_521[1:0]) begin
          match_flag_521 = 1'b1;
          addr[521] = loop_521[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_522 = 1'b0;
        addr[522] = 3'b0;
        for (loop_522 = 0; loop_522 < NUM_CELL; loop_522++) begin
         if ({b[10],a[16]}) == loop_522[1:0]) begin
          match_flag_522 = 1'b1;
          addr[522] = loop_522[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_523 = 1'b0;
        addr[523] = 3'b0;
        for (loop_523 = 0; loop_523 < NUM_CELL; loop_523++) begin
         if ({b[11],a[16]}) == loop_523[1:0]) begin
          match_flag_523 = 1'b1;
          addr[523] = loop_523[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_524 = 1'b0;
        addr[524] = 3'b0;
        for (loop_524 = 0; loop_524 < NUM_CELL; loop_524++) begin
         if ({b[12],a[16]}) == loop_524[1:0]) begin
          match_flag_524 = 1'b1;
          addr[524] = loop_524[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_525 = 1'b0;
        addr[525] = 3'b0;
        for (loop_525 = 0; loop_525 < NUM_CELL; loop_525++) begin
         if ({b[13],a[16]}) == loop_525[1:0]) begin
          match_flag_525 = 1'b1;
          addr[525] = loop_525[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_526 = 1'b0;
        addr[526] = 3'b0;
        for (loop_526 = 0; loop_526 < NUM_CELL; loop_526++) begin
         if ({b[14],a[16]}) == loop_526[1:0]) begin
          match_flag_526 = 1'b1;
          addr[526] = loop_526[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_527 = 1'b0;
        addr[527] = 3'b0;
        for (loop_527 = 0; loop_527 < NUM_CELL; loop_527++) begin
         if ({b[15],a[16]}) == loop_527[1:0]) begin
          match_flag_527 = 1'b1;
          addr[527] = loop_527[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_528 = 1'b0;
        addr[528] = 3'b0;
        for (loop_528 = 0; loop_528 < NUM_CELL; loop_528++) begin
         if ({b[16],a[16]}) == loop_528[1:0]) begin
          match_flag_528 = 1'b1;
          addr[528] = loop_528[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_529 = 1'b0;
        addr[529] = 3'b0;
        for (loop_529 = 0; loop_529 < NUM_CELL; loop_529++) begin
         if ({b[17],a[16]}) == loop_529[1:0]) begin
          match_flag_529 = 1'b1;
          addr[529] = loop_529[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_530 = 1'b0;
        addr[530] = 3'b0;
        for (loop_530 = 0; loop_530 < NUM_CELL; loop_530++) begin
         if ({b[18],a[16]}) == loop_530[1:0]) begin
          match_flag_530 = 1'b1;
          addr[530] = loop_530[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_531 = 1'b0;
        addr[531] = 3'b0;
        for (loop_531 = 0; loop_531 < NUM_CELL; loop_531++) begin
         if ({b[19],a[16]}) == loop_531[1:0]) begin
          match_flag_531 = 1'b1;
          addr[531] = loop_531[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_532 = 1'b0;
        addr[532] = 3'b0;
        for (loop_532 = 0; loop_532 < NUM_CELL; loop_532++) begin
         if ({b[20],a[16]}) == loop_532[1:0]) begin
          match_flag_532 = 1'b1;
          addr[532] = loop_532[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_533 = 1'b0;
        addr[533] = 3'b0;
        for (loop_533 = 0; loop_533 < NUM_CELL; loop_533++) begin
         if ({b[21],a[16]}) == loop_533[1:0]) begin
          match_flag_533 = 1'b1;
          addr[533] = loop_533[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_534 = 1'b0;
        addr[534] = 3'b0;
        for (loop_534 = 0; loop_534 < NUM_CELL; loop_534++) begin
         if ({b[22],a[16]}) == loop_534[1:0]) begin
          match_flag_534 = 1'b1;
          addr[534] = loop_534[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_535 = 1'b0;
        addr[535] = 3'b0;
        for (loop_535 = 0; loop_535 < NUM_CELL; loop_535++) begin
         if ({b[23],a[16]}) == loop_535[1:0]) begin
          match_flag_535 = 1'b1;
          addr[535] = loop_535[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_536 = 1'b0;
        addr[536] = 3'b0;
        for (loop_536 = 0; loop_536 < NUM_CELL; loop_536++) begin
         if ({b[24],a[16]}) == loop_536[1:0]) begin
          match_flag_536 = 1'b1;
          addr[536] = loop_536[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_537 = 1'b0;
        addr[537] = 3'b0;
        for (loop_537 = 0; loop_537 < NUM_CELL; loop_537++) begin
         if ({b[25],a[16]}) == loop_537[1:0]) begin
          match_flag_537 = 1'b1;
          addr[537] = loop_537[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_538 = 1'b0;
        addr[538] = 3'b0;
        for (loop_538 = 0; loop_538 < NUM_CELL; loop_538++) begin
         if ({b[26],a[16]}) == loop_538[1:0]) begin
          match_flag_538 = 1'b1;
          addr[538] = loop_538[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_539 = 1'b0;
        addr[539] = 3'b0;
        for (loop_539 = 0; loop_539 < NUM_CELL; loop_539++) begin
         if ({b[27],a[16]}) == loop_539[1:0]) begin
          match_flag_539 = 1'b1;
          addr[539] = loop_539[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_540 = 1'b0;
        addr[540] = 3'b0;
        for (loop_540 = 0; loop_540 < NUM_CELL; loop_540++) begin
         if ({b[28],a[16]}) == loop_540[1:0]) begin
          match_flag_540 = 1'b1;
          addr[540] = loop_540[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_541 = 1'b0;
        addr[541] = 3'b0;
        for (loop_541 = 0; loop_541 < NUM_CELL; loop_541++) begin
         if ({b[29],a[16]}) == loop_541[1:0]) begin
          match_flag_541 = 1'b1;
          addr[541] = loop_541[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_542 = 1'b0;
        addr[542] = 3'b0;
        for (loop_542 = 0; loop_542 < NUM_CELL; loop_542++) begin
         if ({b[30],a[16]}) == loop_542[1:0]) begin
          match_flag_542 = 1'b1;
          addr[542] = loop_542[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_543 = 1'b0;
        addr[543] = 3'b0;
        for (loop_543 = 0; loop_543 < NUM_CELL; loop_543++) begin
         if ({b[31],a[16]}) == loop_543[1:0]) begin
          match_flag_543 = 1'b1;
          addr[543] = loop_543[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_544 = 1'b0;
        addr[544] = 3'b0;
        for (loop_544 = 0; loop_544 < NUM_CELL; loop_544++) begin
         if ({b[0],a[17]}) == loop_544[1:0]) begin
          match_flag_544 = 1'b1;
          addr[544] = loop_544[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_545 = 1'b0;
        addr[545] = 3'b0;
        for (loop_545 = 0; loop_545 < NUM_CELL; loop_545++) begin
         if ({b[1],a[17]}) == loop_545[1:0]) begin
          match_flag_545 = 1'b1;
          addr[545] = loop_545[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_546 = 1'b0;
        addr[546] = 3'b0;
        for (loop_546 = 0; loop_546 < NUM_CELL; loop_546++) begin
         if ({b[2],a[17]}) == loop_546[1:0]) begin
          match_flag_546 = 1'b1;
          addr[546] = loop_546[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_547 = 1'b0;
        addr[547] = 3'b0;
        for (loop_547 = 0; loop_547 < NUM_CELL; loop_547++) begin
         if ({b[3],a[17]}) == loop_547[1:0]) begin
          match_flag_547 = 1'b1;
          addr[547] = loop_547[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_548 = 1'b0;
        addr[548] = 3'b0;
        for (loop_548 = 0; loop_548 < NUM_CELL; loop_548++) begin
         if ({b[4],a[17]}) == loop_548[1:0]) begin
          match_flag_548 = 1'b1;
          addr[548] = loop_548[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_549 = 1'b0;
        addr[549] = 3'b0;
        for (loop_549 = 0; loop_549 < NUM_CELL; loop_549++) begin
         if ({b[5],a[17]}) == loop_549[1:0]) begin
          match_flag_549 = 1'b1;
          addr[549] = loop_549[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_550 = 1'b0;
        addr[550] = 3'b0;
        for (loop_550 = 0; loop_550 < NUM_CELL; loop_550++) begin
         if ({b[6],a[17]}) == loop_550[1:0]) begin
          match_flag_550 = 1'b1;
          addr[550] = loop_550[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_551 = 1'b0;
        addr[551] = 3'b0;
        for (loop_551 = 0; loop_551 < NUM_CELL; loop_551++) begin
         if ({b[7],a[17]}) == loop_551[1:0]) begin
          match_flag_551 = 1'b1;
          addr[551] = loop_551[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_552 = 1'b0;
        addr[552] = 3'b0;
        for (loop_552 = 0; loop_552 < NUM_CELL; loop_552++) begin
         if ({b[8],a[17]}) == loop_552[1:0]) begin
          match_flag_552 = 1'b1;
          addr[552] = loop_552[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_553 = 1'b0;
        addr[553] = 3'b0;
        for (loop_553 = 0; loop_553 < NUM_CELL; loop_553++) begin
         if ({b[9],a[17]}) == loop_553[1:0]) begin
          match_flag_553 = 1'b1;
          addr[553] = loop_553[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_554 = 1'b0;
        addr[554] = 3'b0;
        for (loop_554 = 0; loop_554 < NUM_CELL; loop_554++) begin
         if ({b[10],a[17]}) == loop_554[1:0]) begin
          match_flag_554 = 1'b1;
          addr[554] = loop_554[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_555 = 1'b0;
        addr[555] = 3'b0;
        for (loop_555 = 0; loop_555 < NUM_CELL; loop_555++) begin
         if ({b[11],a[17]}) == loop_555[1:0]) begin
          match_flag_555 = 1'b1;
          addr[555] = loop_555[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_556 = 1'b0;
        addr[556] = 3'b0;
        for (loop_556 = 0; loop_556 < NUM_CELL; loop_556++) begin
         if ({b[12],a[17]}) == loop_556[1:0]) begin
          match_flag_556 = 1'b1;
          addr[556] = loop_556[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_557 = 1'b0;
        addr[557] = 3'b0;
        for (loop_557 = 0; loop_557 < NUM_CELL; loop_557++) begin
         if ({b[13],a[17]}) == loop_557[1:0]) begin
          match_flag_557 = 1'b1;
          addr[557] = loop_557[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_558 = 1'b0;
        addr[558] = 3'b0;
        for (loop_558 = 0; loop_558 < NUM_CELL; loop_558++) begin
         if ({b[14],a[17]}) == loop_558[1:0]) begin
          match_flag_558 = 1'b1;
          addr[558] = loop_558[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_559 = 1'b0;
        addr[559] = 3'b0;
        for (loop_559 = 0; loop_559 < NUM_CELL; loop_559++) begin
         if ({b[15],a[17]}) == loop_559[1:0]) begin
          match_flag_559 = 1'b1;
          addr[559] = loop_559[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_560 = 1'b0;
        addr[560] = 3'b0;
        for (loop_560 = 0; loop_560 < NUM_CELL; loop_560++) begin
         if ({b[16],a[17]}) == loop_560[1:0]) begin
          match_flag_560 = 1'b1;
          addr[560] = loop_560[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_561 = 1'b0;
        addr[561] = 3'b0;
        for (loop_561 = 0; loop_561 < NUM_CELL; loop_561++) begin
         if ({b[17],a[17]}) == loop_561[1:0]) begin
          match_flag_561 = 1'b1;
          addr[561] = loop_561[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_562 = 1'b0;
        addr[562] = 3'b0;
        for (loop_562 = 0; loop_562 < NUM_CELL; loop_562++) begin
         if ({b[18],a[17]}) == loop_562[1:0]) begin
          match_flag_562 = 1'b1;
          addr[562] = loop_562[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_563 = 1'b0;
        addr[563] = 3'b0;
        for (loop_563 = 0; loop_563 < NUM_CELL; loop_563++) begin
         if ({b[19],a[17]}) == loop_563[1:0]) begin
          match_flag_563 = 1'b1;
          addr[563] = loop_563[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_564 = 1'b0;
        addr[564] = 3'b0;
        for (loop_564 = 0; loop_564 < NUM_CELL; loop_564++) begin
         if ({b[20],a[17]}) == loop_564[1:0]) begin
          match_flag_564 = 1'b1;
          addr[564] = loop_564[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_565 = 1'b0;
        addr[565] = 3'b0;
        for (loop_565 = 0; loop_565 < NUM_CELL; loop_565++) begin
         if ({b[21],a[17]}) == loop_565[1:0]) begin
          match_flag_565 = 1'b1;
          addr[565] = loop_565[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_566 = 1'b0;
        addr[566] = 3'b0;
        for (loop_566 = 0; loop_566 < NUM_CELL; loop_566++) begin
         if ({b[22],a[17]}) == loop_566[1:0]) begin
          match_flag_566 = 1'b1;
          addr[566] = loop_566[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_567 = 1'b0;
        addr[567] = 3'b0;
        for (loop_567 = 0; loop_567 < NUM_CELL; loop_567++) begin
         if ({b[23],a[17]}) == loop_567[1:0]) begin
          match_flag_567 = 1'b1;
          addr[567] = loop_567[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_568 = 1'b0;
        addr[568] = 3'b0;
        for (loop_568 = 0; loop_568 < NUM_CELL; loop_568++) begin
         if ({b[24],a[17]}) == loop_568[1:0]) begin
          match_flag_568 = 1'b1;
          addr[568] = loop_568[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_569 = 1'b0;
        addr[569] = 3'b0;
        for (loop_569 = 0; loop_569 < NUM_CELL; loop_569++) begin
         if ({b[25],a[17]}) == loop_569[1:0]) begin
          match_flag_569 = 1'b1;
          addr[569] = loop_569[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_570 = 1'b0;
        addr[570] = 3'b0;
        for (loop_570 = 0; loop_570 < NUM_CELL; loop_570++) begin
         if ({b[26],a[17]}) == loop_570[1:0]) begin
          match_flag_570 = 1'b1;
          addr[570] = loop_570[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_571 = 1'b0;
        addr[571] = 3'b0;
        for (loop_571 = 0; loop_571 < NUM_CELL; loop_571++) begin
         if ({b[27],a[17]}) == loop_571[1:0]) begin
          match_flag_571 = 1'b1;
          addr[571] = loop_571[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_572 = 1'b0;
        addr[572] = 3'b0;
        for (loop_572 = 0; loop_572 < NUM_CELL; loop_572++) begin
         if ({b[28],a[17]}) == loop_572[1:0]) begin
          match_flag_572 = 1'b1;
          addr[572] = loop_572[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_573 = 1'b0;
        addr[573] = 3'b0;
        for (loop_573 = 0; loop_573 < NUM_CELL; loop_573++) begin
         if ({b[29],a[17]}) == loop_573[1:0]) begin
          match_flag_573 = 1'b1;
          addr[573] = loop_573[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_574 = 1'b0;
        addr[574] = 3'b0;
        for (loop_574 = 0; loop_574 < NUM_CELL; loop_574++) begin
         if ({b[30],a[17]}) == loop_574[1:0]) begin
          match_flag_574 = 1'b1;
          addr[574] = loop_574[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_575 = 1'b0;
        addr[575] = 3'b0;
        for (loop_575 = 0; loop_575 < NUM_CELL; loop_575++) begin
         if ({b[31],a[17]}) == loop_575[1:0]) begin
          match_flag_575 = 1'b1;
          addr[575] = loop_575[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_576 = 1'b0;
        addr[576] = 3'b0;
        for (loop_576 = 0; loop_576 < NUM_CELL; loop_576++) begin
         if ({b[0],a[18]}) == loop_576[1:0]) begin
          match_flag_576 = 1'b1;
          addr[576] = loop_576[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_577 = 1'b0;
        addr[577] = 3'b0;
        for (loop_577 = 0; loop_577 < NUM_CELL; loop_577++) begin
         if ({b[1],a[18]}) == loop_577[1:0]) begin
          match_flag_577 = 1'b1;
          addr[577] = loop_577[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_578 = 1'b0;
        addr[578] = 3'b0;
        for (loop_578 = 0; loop_578 < NUM_CELL; loop_578++) begin
         if ({b[2],a[18]}) == loop_578[1:0]) begin
          match_flag_578 = 1'b1;
          addr[578] = loop_578[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_579 = 1'b0;
        addr[579] = 3'b0;
        for (loop_579 = 0; loop_579 < NUM_CELL; loop_579++) begin
         if ({b[3],a[18]}) == loop_579[1:0]) begin
          match_flag_579 = 1'b1;
          addr[579] = loop_579[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_580 = 1'b0;
        addr[580] = 3'b0;
        for (loop_580 = 0; loop_580 < NUM_CELL; loop_580++) begin
         if ({b[4],a[18]}) == loop_580[1:0]) begin
          match_flag_580 = 1'b1;
          addr[580] = loop_580[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_581 = 1'b0;
        addr[581] = 3'b0;
        for (loop_581 = 0; loop_581 < NUM_CELL; loop_581++) begin
         if ({b[5],a[18]}) == loop_581[1:0]) begin
          match_flag_581 = 1'b1;
          addr[581] = loop_581[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_582 = 1'b0;
        addr[582] = 3'b0;
        for (loop_582 = 0; loop_582 < NUM_CELL; loop_582++) begin
         if ({b[6],a[18]}) == loop_582[1:0]) begin
          match_flag_582 = 1'b1;
          addr[582] = loop_582[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_583 = 1'b0;
        addr[583] = 3'b0;
        for (loop_583 = 0; loop_583 < NUM_CELL; loop_583++) begin
         if ({b[7],a[18]}) == loop_583[1:0]) begin
          match_flag_583 = 1'b1;
          addr[583] = loop_583[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_584 = 1'b0;
        addr[584] = 3'b0;
        for (loop_584 = 0; loop_584 < NUM_CELL; loop_584++) begin
         if ({b[8],a[18]}) == loop_584[1:0]) begin
          match_flag_584 = 1'b1;
          addr[584] = loop_584[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_585 = 1'b0;
        addr[585] = 3'b0;
        for (loop_585 = 0; loop_585 < NUM_CELL; loop_585++) begin
         if ({b[9],a[18]}) == loop_585[1:0]) begin
          match_flag_585 = 1'b1;
          addr[585] = loop_585[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_586 = 1'b0;
        addr[586] = 3'b0;
        for (loop_586 = 0; loop_586 < NUM_CELL; loop_586++) begin
         if ({b[10],a[18]}) == loop_586[1:0]) begin
          match_flag_586 = 1'b1;
          addr[586] = loop_586[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_587 = 1'b0;
        addr[587] = 3'b0;
        for (loop_587 = 0; loop_587 < NUM_CELL; loop_587++) begin
         if ({b[11],a[18]}) == loop_587[1:0]) begin
          match_flag_587 = 1'b1;
          addr[587] = loop_587[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_588 = 1'b0;
        addr[588] = 3'b0;
        for (loop_588 = 0; loop_588 < NUM_CELL; loop_588++) begin
         if ({b[12],a[18]}) == loop_588[1:0]) begin
          match_flag_588 = 1'b1;
          addr[588] = loop_588[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_589 = 1'b0;
        addr[589] = 3'b0;
        for (loop_589 = 0; loop_589 < NUM_CELL; loop_589++) begin
         if ({b[13],a[18]}) == loop_589[1:0]) begin
          match_flag_589 = 1'b1;
          addr[589] = loop_589[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_590 = 1'b0;
        addr[590] = 3'b0;
        for (loop_590 = 0; loop_590 < NUM_CELL; loop_590++) begin
         if ({b[14],a[18]}) == loop_590[1:0]) begin
          match_flag_590 = 1'b1;
          addr[590] = loop_590[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_591 = 1'b0;
        addr[591] = 3'b0;
        for (loop_591 = 0; loop_591 < NUM_CELL; loop_591++) begin
         if ({b[15],a[18]}) == loop_591[1:0]) begin
          match_flag_591 = 1'b1;
          addr[591] = loop_591[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_592 = 1'b0;
        addr[592] = 3'b0;
        for (loop_592 = 0; loop_592 < NUM_CELL; loop_592++) begin
         if ({b[16],a[18]}) == loop_592[1:0]) begin
          match_flag_592 = 1'b1;
          addr[592] = loop_592[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_593 = 1'b0;
        addr[593] = 3'b0;
        for (loop_593 = 0; loop_593 < NUM_CELL; loop_593++) begin
         if ({b[17],a[18]}) == loop_593[1:0]) begin
          match_flag_593 = 1'b1;
          addr[593] = loop_593[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_594 = 1'b0;
        addr[594] = 3'b0;
        for (loop_594 = 0; loop_594 < NUM_CELL; loop_594++) begin
         if ({b[18],a[18]}) == loop_594[1:0]) begin
          match_flag_594 = 1'b1;
          addr[594] = loop_594[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_595 = 1'b0;
        addr[595] = 3'b0;
        for (loop_595 = 0; loop_595 < NUM_CELL; loop_595++) begin
         if ({b[19],a[18]}) == loop_595[1:0]) begin
          match_flag_595 = 1'b1;
          addr[595] = loop_595[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_596 = 1'b0;
        addr[596] = 3'b0;
        for (loop_596 = 0; loop_596 < NUM_CELL; loop_596++) begin
         if ({b[20],a[18]}) == loop_596[1:0]) begin
          match_flag_596 = 1'b1;
          addr[596] = loop_596[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_597 = 1'b0;
        addr[597] = 3'b0;
        for (loop_597 = 0; loop_597 < NUM_CELL; loop_597++) begin
         if ({b[21],a[18]}) == loop_597[1:0]) begin
          match_flag_597 = 1'b1;
          addr[597] = loop_597[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_598 = 1'b0;
        addr[598] = 3'b0;
        for (loop_598 = 0; loop_598 < NUM_CELL; loop_598++) begin
         if ({b[22],a[18]}) == loop_598[1:0]) begin
          match_flag_598 = 1'b1;
          addr[598] = loop_598[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_599 = 1'b0;
        addr[599] = 3'b0;
        for (loop_599 = 0; loop_599 < NUM_CELL; loop_599++) begin
         if ({b[23],a[18]}) == loop_599[1:0]) begin
          match_flag_599 = 1'b1;
          addr[599] = loop_599[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_600 = 1'b0;
        addr[600] = 3'b0;
        for (loop_600 = 0; loop_600 < NUM_CELL; loop_600++) begin
         if ({b[24],a[18]}) == loop_600[1:0]) begin
          match_flag_600 = 1'b1;
          addr[600] = loop_600[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_601 = 1'b0;
        addr[601] = 3'b0;
        for (loop_601 = 0; loop_601 < NUM_CELL; loop_601++) begin
         if ({b[25],a[18]}) == loop_601[1:0]) begin
          match_flag_601 = 1'b1;
          addr[601] = loop_601[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_602 = 1'b0;
        addr[602] = 3'b0;
        for (loop_602 = 0; loop_602 < NUM_CELL; loop_602++) begin
         if ({b[26],a[18]}) == loop_602[1:0]) begin
          match_flag_602 = 1'b1;
          addr[602] = loop_602[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_603 = 1'b0;
        addr[603] = 3'b0;
        for (loop_603 = 0; loop_603 < NUM_CELL; loop_603++) begin
         if ({b[27],a[18]}) == loop_603[1:0]) begin
          match_flag_603 = 1'b1;
          addr[603] = loop_603[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_604 = 1'b0;
        addr[604] = 3'b0;
        for (loop_604 = 0; loop_604 < NUM_CELL; loop_604++) begin
         if ({b[28],a[18]}) == loop_604[1:0]) begin
          match_flag_604 = 1'b1;
          addr[604] = loop_604[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_605 = 1'b0;
        addr[605] = 3'b0;
        for (loop_605 = 0; loop_605 < NUM_CELL; loop_605++) begin
         if ({b[29],a[18]}) == loop_605[1:0]) begin
          match_flag_605 = 1'b1;
          addr[605] = loop_605[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_606 = 1'b0;
        addr[606] = 3'b0;
        for (loop_606 = 0; loop_606 < NUM_CELL; loop_606++) begin
         if ({b[30],a[18]}) == loop_606[1:0]) begin
          match_flag_606 = 1'b1;
          addr[606] = loop_606[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_607 = 1'b0;
        addr[607] = 3'b0;
        for (loop_607 = 0; loop_607 < NUM_CELL; loop_607++) begin
         if ({b[31],a[18]}) == loop_607[1:0]) begin
          match_flag_607 = 1'b1;
          addr[607] = loop_607[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_608 = 1'b0;
        addr[608] = 3'b0;
        for (loop_608 = 0; loop_608 < NUM_CELL; loop_608++) begin
         if ({b[0],a[19]}) == loop_608[1:0]) begin
          match_flag_608 = 1'b1;
          addr[608] = loop_608[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_609 = 1'b0;
        addr[609] = 3'b0;
        for (loop_609 = 0; loop_609 < NUM_CELL; loop_609++) begin
         if ({b[1],a[19]}) == loop_609[1:0]) begin
          match_flag_609 = 1'b1;
          addr[609] = loop_609[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_610 = 1'b0;
        addr[610] = 3'b0;
        for (loop_610 = 0; loop_610 < NUM_CELL; loop_610++) begin
         if ({b[2],a[19]}) == loop_610[1:0]) begin
          match_flag_610 = 1'b1;
          addr[610] = loop_610[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_611 = 1'b0;
        addr[611] = 3'b0;
        for (loop_611 = 0; loop_611 < NUM_CELL; loop_611++) begin
         if ({b[3],a[19]}) == loop_611[1:0]) begin
          match_flag_611 = 1'b1;
          addr[611] = loop_611[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_612 = 1'b0;
        addr[612] = 3'b0;
        for (loop_612 = 0; loop_612 < NUM_CELL; loop_612++) begin
         if ({b[4],a[19]}) == loop_612[1:0]) begin
          match_flag_612 = 1'b1;
          addr[612] = loop_612[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_613 = 1'b0;
        addr[613] = 3'b0;
        for (loop_613 = 0; loop_613 < NUM_CELL; loop_613++) begin
         if ({b[5],a[19]}) == loop_613[1:0]) begin
          match_flag_613 = 1'b1;
          addr[613] = loop_613[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_614 = 1'b0;
        addr[614] = 3'b0;
        for (loop_614 = 0; loop_614 < NUM_CELL; loop_614++) begin
         if ({b[6],a[19]}) == loop_614[1:0]) begin
          match_flag_614 = 1'b1;
          addr[614] = loop_614[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_615 = 1'b0;
        addr[615] = 3'b0;
        for (loop_615 = 0; loop_615 < NUM_CELL; loop_615++) begin
         if ({b[7],a[19]}) == loop_615[1:0]) begin
          match_flag_615 = 1'b1;
          addr[615] = loop_615[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_616 = 1'b0;
        addr[616] = 3'b0;
        for (loop_616 = 0; loop_616 < NUM_CELL; loop_616++) begin
         if ({b[8],a[19]}) == loop_616[1:0]) begin
          match_flag_616 = 1'b1;
          addr[616] = loop_616[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_617 = 1'b0;
        addr[617] = 3'b0;
        for (loop_617 = 0; loop_617 < NUM_CELL; loop_617++) begin
         if ({b[9],a[19]}) == loop_617[1:0]) begin
          match_flag_617 = 1'b1;
          addr[617] = loop_617[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_618 = 1'b0;
        addr[618] = 3'b0;
        for (loop_618 = 0; loop_618 < NUM_CELL; loop_618++) begin
         if ({b[10],a[19]}) == loop_618[1:0]) begin
          match_flag_618 = 1'b1;
          addr[618] = loop_618[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_619 = 1'b0;
        addr[619] = 3'b0;
        for (loop_619 = 0; loop_619 < NUM_CELL; loop_619++) begin
         if ({b[11],a[19]}) == loop_619[1:0]) begin
          match_flag_619 = 1'b1;
          addr[619] = loop_619[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_620 = 1'b0;
        addr[620] = 3'b0;
        for (loop_620 = 0; loop_620 < NUM_CELL; loop_620++) begin
         if ({b[12],a[19]}) == loop_620[1:0]) begin
          match_flag_620 = 1'b1;
          addr[620] = loop_620[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_621 = 1'b0;
        addr[621] = 3'b0;
        for (loop_621 = 0; loop_621 < NUM_CELL; loop_621++) begin
         if ({b[13],a[19]}) == loop_621[1:0]) begin
          match_flag_621 = 1'b1;
          addr[621] = loop_621[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_622 = 1'b0;
        addr[622] = 3'b0;
        for (loop_622 = 0; loop_622 < NUM_CELL; loop_622++) begin
         if ({b[14],a[19]}) == loop_622[1:0]) begin
          match_flag_622 = 1'b1;
          addr[622] = loop_622[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_623 = 1'b0;
        addr[623] = 3'b0;
        for (loop_623 = 0; loop_623 < NUM_CELL; loop_623++) begin
         if ({b[15],a[19]}) == loop_623[1:0]) begin
          match_flag_623 = 1'b1;
          addr[623] = loop_623[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_624 = 1'b0;
        addr[624] = 3'b0;
        for (loop_624 = 0; loop_624 < NUM_CELL; loop_624++) begin
         if ({b[16],a[19]}) == loop_624[1:0]) begin
          match_flag_624 = 1'b1;
          addr[624] = loop_624[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_625 = 1'b0;
        addr[625] = 3'b0;
        for (loop_625 = 0; loop_625 < NUM_CELL; loop_625++) begin
         if ({b[17],a[19]}) == loop_625[1:0]) begin
          match_flag_625 = 1'b1;
          addr[625] = loop_625[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_626 = 1'b0;
        addr[626] = 3'b0;
        for (loop_626 = 0; loop_626 < NUM_CELL; loop_626++) begin
         if ({b[18],a[19]}) == loop_626[1:0]) begin
          match_flag_626 = 1'b1;
          addr[626] = loop_626[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_627 = 1'b0;
        addr[627] = 3'b0;
        for (loop_627 = 0; loop_627 < NUM_CELL; loop_627++) begin
         if ({b[19],a[19]}) == loop_627[1:0]) begin
          match_flag_627 = 1'b1;
          addr[627] = loop_627[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_628 = 1'b0;
        addr[628] = 3'b0;
        for (loop_628 = 0; loop_628 < NUM_CELL; loop_628++) begin
         if ({b[20],a[19]}) == loop_628[1:0]) begin
          match_flag_628 = 1'b1;
          addr[628] = loop_628[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_629 = 1'b0;
        addr[629] = 3'b0;
        for (loop_629 = 0; loop_629 < NUM_CELL; loop_629++) begin
         if ({b[21],a[19]}) == loop_629[1:0]) begin
          match_flag_629 = 1'b1;
          addr[629] = loop_629[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_630 = 1'b0;
        addr[630] = 3'b0;
        for (loop_630 = 0; loop_630 < NUM_CELL; loop_630++) begin
         if ({b[22],a[19]}) == loop_630[1:0]) begin
          match_flag_630 = 1'b1;
          addr[630] = loop_630[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_631 = 1'b0;
        addr[631] = 3'b0;
        for (loop_631 = 0; loop_631 < NUM_CELL; loop_631++) begin
         if ({b[23],a[19]}) == loop_631[1:0]) begin
          match_flag_631 = 1'b1;
          addr[631] = loop_631[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_632 = 1'b0;
        addr[632] = 3'b0;
        for (loop_632 = 0; loop_632 < NUM_CELL; loop_632++) begin
         if ({b[24],a[19]}) == loop_632[1:0]) begin
          match_flag_632 = 1'b1;
          addr[632] = loop_632[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_633 = 1'b0;
        addr[633] = 3'b0;
        for (loop_633 = 0; loop_633 < NUM_CELL; loop_633++) begin
         if ({b[25],a[19]}) == loop_633[1:0]) begin
          match_flag_633 = 1'b1;
          addr[633] = loop_633[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_634 = 1'b0;
        addr[634] = 3'b0;
        for (loop_634 = 0; loop_634 < NUM_CELL; loop_634++) begin
         if ({b[26],a[19]}) == loop_634[1:0]) begin
          match_flag_634 = 1'b1;
          addr[634] = loop_634[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_635 = 1'b0;
        addr[635] = 3'b0;
        for (loop_635 = 0; loop_635 < NUM_CELL; loop_635++) begin
         if ({b[27],a[19]}) == loop_635[1:0]) begin
          match_flag_635 = 1'b1;
          addr[635] = loop_635[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_636 = 1'b0;
        addr[636] = 3'b0;
        for (loop_636 = 0; loop_636 < NUM_CELL; loop_636++) begin
         if ({b[28],a[19]}) == loop_636[1:0]) begin
          match_flag_636 = 1'b1;
          addr[636] = loop_636[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_637 = 1'b0;
        addr[637] = 3'b0;
        for (loop_637 = 0; loop_637 < NUM_CELL; loop_637++) begin
         if ({b[29],a[19]}) == loop_637[1:0]) begin
          match_flag_637 = 1'b1;
          addr[637] = loop_637[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_638 = 1'b0;
        addr[638] = 3'b0;
        for (loop_638 = 0; loop_638 < NUM_CELL; loop_638++) begin
         if ({b[30],a[19]}) == loop_638[1:0]) begin
          match_flag_638 = 1'b1;
          addr[638] = loop_638[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_639 = 1'b0;
        addr[639] = 3'b0;
        for (loop_639 = 0; loop_639 < NUM_CELL; loop_639++) begin
         if ({b[31],a[19]}) == loop_639[1:0]) begin
          match_flag_639 = 1'b1;
          addr[639] = loop_639[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_640 = 1'b0;
        addr[640] = 3'b0;
        for (loop_640 = 0; loop_640 < NUM_CELL; loop_640++) begin
         if ({b[0],a[20]}) == loop_640[1:0]) begin
          match_flag_640 = 1'b1;
          addr[640] = loop_640[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_641 = 1'b0;
        addr[641] = 3'b0;
        for (loop_641 = 0; loop_641 < NUM_CELL; loop_641++) begin
         if ({b[1],a[20]}) == loop_641[1:0]) begin
          match_flag_641 = 1'b1;
          addr[641] = loop_641[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_642 = 1'b0;
        addr[642] = 3'b0;
        for (loop_642 = 0; loop_642 < NUM_CELL; loop_642++) begin
         if ({b[2],a[20]}) == loop_642[1:0]) begin
          match_flag_642 = 1'b1;
          addr[642] = loop_642[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_643 = 1'b0;
        addr[643] = 3'b0;
        for (loop_643 = 0; loop_643 < NUM_CELL; loop_643++) begin
         if ({b[3],a[20]}) == loop_643[1:0]) begin
          match_flag_643 = 1'b1;
          addr[643] = loop_643[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_644 = 1'b0;
        addr[644] = 3'b0;
        for (loop_644 = 0; loop_644 < NUM_CELL; loop_644++) begin
         if ({b[4],a[20]}) == loop_644[1:0]) begin
          match_flag_644 = 1'b1;
          addr[644] = loop_644[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_645 = 1'b0;
        addr[645] = 3'b0;
        for (loop_645 = 0; loop_645 < NUM_CELL; loop_645++) begin
         if ({b[5],a[20]}) == loop_645[1:0]) begin
          match_flag_645 = 1'b1;
          addr[645] = loop_645[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_646 = 1'b0;
        addr[646] = 3'b0;
        for (loop_646 = 0; loop_646 < NUM_CELL; loop_646++) begin
         if ({b[6],a[20]}) == loop_646[1:0]) begin
          match_flag_646 = 1'b1;
          addr[646] = loop_646[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_647 = 1'b0;
        addr[647] = 3'b0;
        for (loop_647 = 0; loop_647 < NUM_CELL; loop_647++) begin
         if ({b[7],a[20]}) == loop_647[1:0]) begin
          match_flag_647 = 1'b1;
          addr[647] = loop_647[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_648 = 1'b0;
        addr[648] = 3'b0;
        for (loop_648 = 0; loop_648 < NUM_CELL; loop_648++) begin
         if ({b[8],a[20]}) == loop_648[1:0]) begin
          match_flag_648 = 1'b1;
          addr[648] = loop_648[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_649 = 1'b0;
        addr[649] = 3'b0;
        for (loop_649 = 0; loop_649 < NUM_CELL; loop_649++) begin
         if ({b[9],a[20]}) == loop_649[1:0]) begin
          match_flag_649 = 1'b1;
          addr[649] = loop_649[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_650 = 1'b0;
        addr[650] = 3'b0;
        for (loop_650 = 0; loop_650 < NUM_CELL; loop_650++) begin
         if ({b[10],a[20]}) == loop_650[1:0]) begin
          match_flag_650 = 1'b1;
          addr[650] = loop_650[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_651 = 1'b0;
        addr[651] = 3'b0;
        for (loop_651 = 0; loop_651 < NUM_CELL; loop_651++) begin
         if ({b[11],a[20]}) == loop_651[1:0]) begin
          match_flag_651 = 1'b1;
          addr[651] = loop_651[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_652 = 1'b0;
        addr[652] = 3'b0;
        for (loop_652 = 0; loop_652 < NUM_CELL; loop_652++) begin
         if ({b[12],a[20]}) == loop_652[1:0]) begin
          match_flag_652 = 1'b1;
          addr[652] = loop_652[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_653 = 1'b0;
        addr[653] = 3'b0;
        for (loop_653 = 0; loop_653 < NUM_CELL; loop_653++) begin
         if ({b[13],a[20]}) == loop_653[1:0]) begin
          match_flag_653 = 1'b1;
          addr[653] = loop_653[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_654 = 1'b0;
        addr[654] = 3'b0;
        for (loop_654 = 0; loop_654 < NUM_CELL; loop_654++) begin
         if ({b[14],a[20]}) == loop_654[1:0]) begin
          match_flag_654 = 1'b1;
          addr[654] = loop_654[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_655 = 1'b0;
        addr[655] = 3'b0;
        for (loop_655 = 0; loop_655 < NUM_CELL; loop_655++) begin
         if ({b[15],a[20]}) == loop_655[1:0]) begin
          match_flag_655 = 1'b1;
          addr[655] = loop_655[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_656 = 1'b0;
        addr[656] = 3'b0;
        for (loop_656 = 0; loop_656 < NUM_CELL; loop_656++) begin
         if ({b[16],a[20]}) == loop_656[1:0]) begin
          match_flag_656 = 1'b1;
          addr[656] = loop_656[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_657 = 1'b0;
        addr[657] = 3'b0;
        for (loop_657 = 0; loop_657 < NUM_CELL; loop_657++) begin
         if ({b[17],a[20]}) == loop_657[1:0]) begin
          match_flag_657 = 1'b1;
          addr[657] = loop_657[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_658 = 1'b0;
        addr[658] = 3'b0;
        for (loop_658 = 0; loop_658 < NUM_CELL; loop_658++) begin
         if ({b[18],a[20]}) == loop_658[1:0]) begin
          match_flag_658 = 1'b1;
          addr[658] = loop_658[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_659 = 1'b0;
        addr[659] = 3'b0;
        for (loop_659 = 0; loop_659 < NUM_CELL; loop_659++) begin
         if ({b[19],a[20]}) == loop_659[1:0]) begin
          match_flag_659 = 1'b1;
          addr[659] = loop_659[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_660 = 1'b0;
        addr[660] = 3'b0;
        for (loop_660 = 0; loop_660 < NUM_CELL; loop_660++) begin
         if ({b[20],a[20]}) == loop_660[1:0]) begin
          match_flag_660 = 1'b1;
          addr[660] = loop_660[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_661 = 1'b0;
        addr[661] = 3'b0;
        for (loop_661 = 0; loop_661 < NUM_CELL; loop_661++) begin
         if ({b[21],a[20]}) == loop_661[1:0]) begin
          match_flag_661 = 1'b1;
          addr[661] = loop_661[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_662 = 1'b0;
        addr[662] = 3'b0;
        for (loop_662 = 0; loop_662 < NUM_CELL; loop_662++) begin
         if ({b[22],a[20]}) == loop_662[1:0]) begin
          match_flag_662 = 1'b1;
          addr[662] = loop_662[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_663 = 1'b0;
        addr[663] = 3'b0;
        for (loop_663 = 0; loop_663 < NUM_CELL; loop_663++) begin
         if ({b[23],a[20]}) == loop_663[1:0]) begin
          match_flag_663 = 1'b1;
          addr[663] = loop_663[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_664 = 1'b0;
        addr[664] = 3'b0;
        for (loop_664 = 0; loop_664 < NUM_CELL; loop_664++) begin
         if ({b[24],a[20]}) == loop_664[1:0]) begin
          match_flag_664 = 1'b1;
          addr[664] = loop_664[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_665 = 1'b0;
        addr[665] = 3'b0;
        for (loop_665 = 0; loop_665 < NUM_CELL; loop_665++) begin
         if ({b[25],a[20]}) == loop_665[1:0]) begin
          match_flag_665 = 1'b1;
          addr[665] = loop_665[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_666 = 1'b0;
        addr[666] = 3'b0;
        for (loop_666 = 0; loop_666 < NUM_CELL; loop_666++) begin
         if ({b[26],a[20]}) == loop_666[1:0]) begin
          match_flag_666 = 1'b1;
          addr[666] = loop_666[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_667 = 1'b0;
        addr[667] = 3'b0;
        for (loop_667 = 0; loop_667 < NUM_CELL; loop_667++) begin
         if ({b[27],a[20]}) == loop_667[1:0]) begin
          match_flag_667 = 1'b1;
          addr[667] = loop_667[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_668 = 1'b0;
        addr[668] = 3'b0;
        for (loop_668 = 0; loop_668 < NUM_CELL; loop_668++) begin
         if ({b[28],a[20]}) == loop_668[1:0]) begin
          match_flag_668 = 1'b1;
          addr[668] = loop_668[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_669 = 1'b0;
        addr[669] = 3'b0;
        for (loop_669 = 0; loop_669 < NUM_CELL; loop_669++) begin
         if ({b[29],a[20]}) == loop_669[1:0]) begin
          match_flag_669 = 1'b1;
          addr[669] = loop_669[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_670 = 1'b0;
        addr[670] = 3'b0;
        for (loop_670 = 0; loop_670 < NUM_CELL; loop_670++) begin
         if ({b[30],a[20]}) == loop_670[1:0]) begin
          match_flag_670 = 1'b1;
          addr[670] = loop_670[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_671 = 1'b0;
        addr[671] = 3'b0;
        for (loop_671 = 0; loop_671 < NUM_CELL; loop_671++) begin
         if ({b[31],a[20]}) == loop_671[1:0]) begin
          match_flag_671 = 1'b1;
          addr[671] = loop_671[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_672 = 1'b0;
        addr[672] = 3'b0;
        for (loop_672 = 0; loop_672 < NUM_CELL; loop_672++) begin
         if ({b[0],a[21]}) == loop_672[1:0]) begin
          match_flag_672 = 1'b1;
          addr[672] = loop_672[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_673 = 1'b0;
        addr[673] = 3'b0;
        for (loop_673 = 0; loop_673 < NUM_CELL; loop_673++) begin
         if ({b[1],a[21]}) == loop_673[1:0]) begin
          match_flag_673 = 1'b1;
          addr[673] = loop_673[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_674 = 1'b0;
        addr[674] = 3'b0;
        for (loop_674 = 0; loop_674 < NUM_CELL; loop_674++) begin
         if ({b[2],a[21]}) == loop_674[1:0]) begin
          match_flag_674 = 1'b1;
          addr[674] = loop_674[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_675 = 1'b0;
        addr[675] = 3'b0;
        for (loop_675 = 0; loop_675 < NUM_CELL; loop_675++) begin
         if ({b[3],a[21]}) == loop_675[1:0]) begin
          match_flag_675 = 1'b1;
          addr[675] = loop_675[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_676 = 1'b0;
        addr[676] = 3'b0;
        for (loop_676 = 0; loop_676 < NUM_CELL; loop_676++) begin
         if ({b[4],a[21]}) == loop_676[1:0]) begin
          match_flag_676 = 1'b1;
          addr[676] = loop_676[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_677 = 1'b0;
        addr[677] = 3'b0;
        for (loop_677 = 0; loop_677 < NUM_CELL; loop_677++) begin
         if ({b[5],a[21]}) == loop_677[1:0]) begin
          match_flag_677 = 1'b1;
          addr[677] = loop_677[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_678 = 1'b0;
        addr[678] = 3'b0;
        for (loop_678 = 0; loop_678 < NUM_CELL; loop_678++) begin
         if ({b[6],a[21]}) == loop_678[1:0]) begin
          match_flag_678 = 1'b1;
          addr[678] = loop_678[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_679 = 1'b0;
        addr[679] = 3'b0;
        for (loop_679 = 0; loop_679 < NUM_CELL; loop_679++) begin
         if ({b[7],a[21]}) == loop_679[1:0]) begin
          match_flag_679 = 1'b1;
          addr[679] = loop_679[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_680 = 1'b0;
        addr[680] = 3'b0;
        for (loop_680 = 0; loop_680 < NUM_CELL; loop_680++) begin
         if ({b[8],a[21]}) == loop_680[1:0]) begin
          match_flag_680 = 1'b1;
          addr[680] = loop_680[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_681 = 1'b0;
        addr[681] = 3'b0;
        for (loop_681 = 0; loop_681 < NUM_CELL; loop_681++) begin
         if ({b[9],a[21]}) == loop_681[1:0]) begin
          match_flag_681 = 1'b1;
          addr[681] = loop_681[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_682 = 1'b0;
        addr[682] = 3'b0;
        for (loop_682 = 0; loop_682 < NUM_CELL; loop_682++) begin
         if ({b[10],a[21]}) == loop_682[1:0]) begin
          match_flag_682 = 1'b1;
          addr[682] = loop_682[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_683 = 1'b0;
        addr[683] = 3'b0;
        for (loop_683 = 0; loop_683 < NUM_CELL; loop_683++) begin
         if ({b[11],a[21]}) == loop_683[1:0]) begin
          match_flag_683 = 1'b1;
          addr[683] = loop_683[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_684 = 1'b0;
        addr[684] = 3'b0;
        for (loop_684 = 0; loop_684 < NUM_CELL; loop_684++) begin
         if ({b[12],a[21]}) == loop_684[1:0]) begin
          match_flag_684 = 1'b1;
          addr[684] = loop_684[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_685 = 1'b0;
        addr[685] = 3'b0;
        for (loop_685 = 0; loop_685 < NUM_CELL; loop_685++) begin
         if ({b[13],a[21]}) == loop_685[1:0]) begin
          match_flag_685 = 1'b1;
          addr[685] = loop_685[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_686 = 1'b0;
        addr[686] = 3'b0;
        for (loop_686 = 0; loop_686 < NUM_CELL; loop_686++) begin
         if ({b[14],a[21]}) == loop_686[1:0]) begin
          match_flag_686 = 1'b1;
          addr[686] = loop_686[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_687 = 1'b0;
        addr[687] = 3'b0;
        for (loop_687 = 0; loop_687 < NUM_CELL; loop_687++) begin
         if ({b[15],a[21]}) == loop_687[1:0]) begin
          match_flag_687 = 1'b1;
          addr[687] = loop_687[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_688 = 1'b0;
        addr[688] = 3'b0;
        for (loop_688 = 0; loop_688 < NUM_CELL; loop_688++) begin
         if ({b[16],a[21]}) == loop_688[1:0]) begin
          match_flag_688 = 1'b1;
          addr[688] = loop_688[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_689 = 1'b0;
        addr[689] = 3'b0;
        for (loop_689 = 0; loop_689 < NUM_CELL; loop_689++) begin
         if ({b[17],a[21]}) == loop_689[1:0]) begin
          match_flag_689 = 1'b1;
          addr[689] = loop_689[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_690 = 1'b0;
        addr[690] = 3'b0;
        for (loop_690 = 0; loop_690 < NUM_CELL; loop_690++) begin
         if ({b[18],a[21]}) == loop_690[1:0]) begin
          match_flag_690 = 1'b1;
          addr[690] = loop_690[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_691 = 1'b0;
        addr[691] = 3'b0;
        for (loop_691 = 0; loop_691 < NUM_CELL; loop_691++) begin
         if ({b[19],a[21]}) == loop_691[1:0]) begin
          match_flag_691 = 1'b1;
          addr[691] = loop_691[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_692 = 1'b0;
        addr[692] = 3'b0;
        for (loop_692 = 0; loop_692 < NUM_CELL; loop_692++) begin
         if ({b[20],a[21]}) == loop_692[1:0]) begin
          match_flag_692 = 1'b1;
          addr[692] = loop_692[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_693 = 1'b0;
        addr[693] = 3'b0;
        for (loop_693 = 0; loop_693 < NUM_CELL; loop_693++) begin
         if ({b[21],a[21]}) == loop_693[1:0]) begin
          match_flag_693 = 1'b1;
          addr[693] = loop_693[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_694 = 1'b0;
        addr[694] = 3'b0;
        for (loop_694 = 0; loop_694 < NUM_CELL; loop_694++) begin
         if ({b[22],a[21]}) == loop_694[1:0]) begin
          match_flag_694 = 1'b1;
          addr[694] = loop_694[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_695 = 1'b0;
        addr[695] = 3'b0;
        for (loop_695 = 0; loop_695 < NUM_CELL; loop_695++) begin
         if ({b[23],a[21]}) == loop_695[1:0]) begin
          match_flag_695 = 1'b1;
          addr[695] = loop_695[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_696 = 1'b0;
        addr[696] = 3'b0;
        for (loop_696 = 0; loop_696 < NUM_CELL; loop_696++) begin
         if ({b[24],a[21]}) == loop_696[1:0]) begin
          match_flag_696 = 1'b1;
          addr[696] = loop_696[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_697 = 1'b0;
        addr[697] = 3'b0;
        for (loop_697 = 0; loop_697 < NUM_CELL; loop_697++) begin
         if ({b[25],a[21]}) == loop_697[1:0]) begin
          match_flag_697 = 1'b1;
          addr[697] = loop_697[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_698 = 1'b0;
        addr[698] = 3'b0;
        for (loop_698 = 0; loop_698 < NUM_CELL; loop_698++) begin
         if ({b[26],a[21]}) == loop_698[1:0]) begin
          match_flag_698 = 1'b1;
          addr[698] = loop_698[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_699 = 1'b0;
        addr[699] = 3'b0;
        for (loop_699 = 0; loop_699 < NUM_CELL; loop_699++) begin
         if ({b[27],a[21]}) == loop_699[1:0]) begin
          match_flag_699 = 1'b1;
          addr[699] = loop_699[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_700 = 1'b0;
        addr[700] = 3'b0;
        for (loop_700 = 0; loop_700 < NUM_CELL; loop_700++) begin
         if ({b[28],a[21]}) == loop_700[1:0]) begin
          match_flag_700 = 1'b1;
          addr[700] = loop_700[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_701 = 1'b0;
        addr[701] = 3'b0;
        for (loop_701 = 0; loop_701 < NUM_CELL; loop_701++) begin
         if ({b[29],a[21]}) == loop_701[1:0]) begin
          match_flag_701 = 1'b1;
          addr[701] = loop_701[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_702 = 1'b0;
        addr[702] = 3'b0;
        for (loop_702 = 0; loop_702 < NUM_CELL; loop_702++) begin
         if ({b[30],a[21]}) == loop_702[1:0]) begin
          match_flag_702 = 1'b1;
          addr[702] = loop_702[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_703 = 1'b0;
        addr[703] = 3'b0;
        for (loop_703 = 0; loop_703 < NUM_CELL; loop_703++) begin
         if ({b[31],a[21]}) == loop_703[1:0]) begin
          match_flag_703 = 1'b1;
          addr[703] = loop_703[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_704 = 1'b0;
        addr[704] = 3'b0;
        for (loop_704 = 0; loop_704 < NUM_CELL; loop_704++) begin
         if ({b[0],a[22]}) == loop_704[1:0]) begin
          match_flag_704 = 1'b1;
          addr[704] = loop_704[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_705 = 1'b0;
        addr[705] = 3'b0;
        for (loop_705 = 0; loop_705 < NUM_CELL; loop_705++) begin
         if ({b[1],a[22]}) == loop_705[1:0]) begin
          match_flag_705 = 1'b1;
          addr[705] = loop_705[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_706 = 1'b0;
        addr[706] = 3'b0;
        for (loop_706 = 0; loop_706 < NUM_CELL; loop_706++) begin
         if ({b[2],a[22]}) == loop_706[1:0]) begin
          match_flag_706 = 1'b1;
          addr[706] = loop_706[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_707 = 1'b0;
        addr[707] = 3'b0;
        for (loop_707 = 0; loop_707 < NUM_CELL; loop_707++) begin
         if ({b[3],a[22]}) == loop_707[1:0]) begin
          match_flag_707 = 1'b1;
          addr[707] = loop_707[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_708 = 1'b0;
        addr[708] = 3'b0;
        for (loop_708 = 0; loop_708 < NUM_CELL; loop_708++) begin
         if ({b[4],a[22]}) == loop_708[1:0]) begin
          match_flag_708 = 1'b1;
          addr[708] = loop_708[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_709 = 1'b0;
        addr[709] = 3'b0;
        for (loop_709 = 0; loop_709 < NUM_CELL; loop_709++) begin
         if ({b[5],a[22]}) == loop_709[1:0]) begin
          match_flag_709 = 1'b1;
          addr[709] = loop_709[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_710 = 1'b0;
        addr[710] = 3'b0;
        for (loop_710 = 0; loop_710 < NUM_CELL; loop_710++) begin
         if ({b[6],a[22]}) == loop_710[1:0]) begin
          match_flag_710 = 1'b1;
          addr[710] = loop_710[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_711 = 1'b0;
        addr[711] = 3'b0;
        for (loop_711 = 0; loop_711 < NUM_CELL; loop_711++) begin
         if ({b[7],a[22]}) == loop_711[1:0]) begin
          match_flag_711 = 1'b1;
          addr[711] = loop_711[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_712 = 1'b0;
        addr[712] = 3'b0;
        for (loop_712 = 0; loop_712 < NUM_CELL; loop_712++) begin
         if ({b[8],a[22]}) == loop_712[1:0]) begin
          match_flag_712 = 1'b1;
          addr[712] = loop_712[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_713 = 1'b0;
        addr[713] = 3'b0;
        for (loop_713 = 0; loop_713 < NUM_CELL; loop_713++) begin
         if ({b[9],a[22]}) == loop_713[1:0]) begin
          match_flag_713 = 1'b1;
          addr[713] = loop_713[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_714 = 1'b0;
        addr[714] = 3'b0;
        for (loop_714 = 0; loop_714 < NUM_CELL; loop_714++) begin
         if ({b[10],a[22]}) == loop_714[1:0]) begin
          match_flag_714 = 1'b1;
          addr[714] = loop_714[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_715 = 1'b0;
        addr[715] = 3'b0;
        for (loop_715 = 0; loop_715 < NUM_CELL; loop_715++) begin
         if ({b[11],a[22]}) == loop_715[1:0]) begin
          match_flag_715 = 1'b1;
          addr[715] = loop_715[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_716 = 1'b0;
        addr[716] = 3'b0;
        for (loop_716 = 0; loop_716 < NUM_CELL; loop_716++) begin
         if ({b[12],a[22]}) == loop_716[1:0]) begin
          match_flag_716 = 1'b1;
          addr[716] = loop_716[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_717 = 1'b0;
        addr[717] = 3'b0;
        for (loop_717 = 0; loop_717 < NUM_CELL; loop_717++) begin
         if ({b[13],a[22]}) == loop_717[1:0]) begin
          match_flag_717 = 1'b1;
          addr[717] = loop_717[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_718 = 1'b0;
        addr[718] = 3'b0;
        for (loop_718 = 0; loop_718 < NUM_CELL; loop_718++) begin
         if ({b[14],a[22]}) == loop_718[1:0]) begin
          match_flag_718 = 1'b1;
          addr[718] = loop_718[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_719 = 1'b0;
        addr[719] = 3'b0;
        for (loop_719 = 0; loop_719 < NUM_CELL; loop_719++) begin
         if ({b[15],a[22]}) == loop_719[1:0]) begin
          match_flag_719 = 1'b1;
          addr[719] = loop_719[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_720 = 1'b0;
        addr[720] = 3'b0;
        for (loop_720 = 0; loop_720 < NUM_CELL; loop_720++) begin
         if ({b[16],a[22]}) == loop_720[1:0]) begin
          match_flag_720 = 1'b1;
          addr[720] = loop_720[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_721 = 1'b0;
        addr[721] = 3'b0;
        for (loop_721 = 0; loop_721 < NUM_CELL; loop_721++) begin
         if ({b[17],a[22]}) == loop_721[1:0]) begin
          match_flag_721 = 1'b1;
          addr[721] = loop_721[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_722 = 1'b0;
        addr[722] = 3'b0;
        for (loop_722 = 0; loop_722 < NUM_CELL; loop_722++) begin
         if ({b[18],a[22]}) == loop_722[1:0]) begin
          match_flag_722 = 1'b1;
          addr[722] = loop_722[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_723 = 1'b0;
        addr[723] = 3'b0;
        for (loop_723 = 0; loop_723 < NUM_CELL; loop_723++) begin
         if ({b[19],a[22]}) == loop_723[1:0]) begin
          match_flag_723 = 1'b1;
          addr[723] = loop_723[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_724 = 1'b0;
        addr[724] = 3'b0;
        for (loop_724 = 0; loop_724 < NUM_CELL; loop_724++) begin
         if ({b[20],a[22]}) == loop_724[1:0]) begin
          match_flag_724 = 1'b1;
          addr[724] = loop_724[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_725 = 1'b0;
        addr[725] = 3'b0;
        for (loop_725 = 0; loop_725 < NUM_CELL; loop_725++) begin
         if ({b[21],a[22]}) == loop_725[1:0]) begin
          match_flag_725 = 1'b1;
          addr[725] = loop_725[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_726 = 1'b0;
        addr[726] = 3'b0;
        for (loop_726 = 0; loop_726 < NUM_CELL; loop_726++) begin
         if ({b[22],a[22]}) == loop_726[1:0]) begin
          match_flag_726 = 1'b1;
          addr[726] = loop_726[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_727 = 1'b0;
        addr[727] = 3'b0;
        for (loop_727 = 0; loop_727 < NUM_CELL; loop_727++) begin
         if ({b[23],a[22]}) == loop_727[1:0]) begin
          match_flag_727 = 1'b1;
          addr[727] = loop_727[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_728 = 1'b0;
        addr[728] = 3'b0;
        for (loop_728 = 0; loop_728 < NUM_CELL; loop_728++) begin
         if ({b[24],a[22]}) == loop_728[1:0]) begin
          match_flag_728 = 1'b1;
          addr[728] = loop_728[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_729 = 1'b0;
        addr[729] = 3'b0;
        for (loop_729 = 0; loop_729 < NUM_CELL; loop_729++) begin
         if ({b[25],a[22]}) == loop_729[1:0]) begin
          match_flag_729 = 1'b1;
          addr[729] = loop_729[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_730 = 1'b0;
        addr[730] = 3'b0;
        for (loop_730 = 0; loop_730 < NUM_CELL; loop_730++) begin
         if ({b[26],a[22]}) == loop_730[1:0]) begin
          match_flag_730 = 1'b1;
          addr[730] = loop_730[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_731 = 1'b0;
        addr[731] = 3'b0;
        for (loop_731 = 0; loop_731 < NUM_CELL; loop_731++) begin
         if ({b[27],a[22]}) == loop_731[1:0]) begin
          match_flag_731 = 1'b1;
          addr[731] = loop_731[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_732 = 1'b0;
        addr[732] = 3'b0;
        for (loop_732 = 0; loop_732 < NUM_CELL; loop_732++) begin
         if ({b[28],a[22]}) == loop_732[1:0]) begin
          match_flag_732 = 1'b1;
          addr[732] = loop_732[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_733 = 1'b0;
        addr[733] = 3'b0;
        for (loop_733 = 0; loop_733 < NUM_CELL; loop_733++) begin
         if ({b[29],a[22]}) == loop_733[1:0]) begin
          match_flag_733 = 1'b1;
          addr[733] = loop_733[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_734 = 1'b0;
        addr[734] = 3'b0;
        for (loop_734 = 0; loop_734 < NUM_CELL; loop_734++) begin
         if ({b[30],a[22]}) == loop_734[1:0]) begin
          match_flag_734 = 1'b1;
          addr[734] = loop_734[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_735 = 1'b0;
        addr[735] = 3'b0;
        for (loop_735 = 0; loop_735 < NUM_CELL; loop_735++) begin
         if ({b[31],a[22]}) == loop_735[1:0]) begin
          match_flag_735 = 1'b1;
          addr[735] = loop_735[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_736 = 1'b0;
        addr[736] = 3'b0;
        for (loop_736 = 0; loop_736 < NUM_CELL; loop_736++) begin
         if ({b[0],a[23]}) == loop_736[1:0]) begin
          match_flag_736 = 1'b1;
          addr[736] = loop_736[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_737 = 1'b0;
        addr[737] = 3'b0;
        for (loop_737 = 0; loop_737 < NUM_CELL; loop_737++) begin
         if ({b[1],a[23]}) == loop_737[1:0]) begin
          match_flag_737 = 1'b1;
          addr[737] = loop_737[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_738 = 1'b0;
        addr[738] = 3'b0;
        for (loop_738 = 0; loop_738 < NUM_CELL; loop_738++) begin
         if ({b[2],a[23]}) == loop_738[1:0]) begin
          match_flag_738 = 1'b1;
          addr[738] = loop_738[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_739 = 1'b0;
        addr[739] = 3'b0;
        for (loop_739 = 0; loop_739 < NUM_CELL; loop_739++) begin
         if ({b[3],a[23]}) == loop_739[1:0]) begin
          match_flag_739 = 1'b1;
          addr[739] = loop_739[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_740 = 1'b0;
        addr[740] = 3'b0;
        for (loop_740 = 0; loop_740 < NUM_CELL; loop_740++) begin
         if ({b[4],a[23]}) == loop_740[1:0]) begin
          match_flag_740 = 1'b1;
          addr[740] = loop_740[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_741 = 1'b0;
        addr[741] = 3'b0;
        for (loop_741 = 0; loop_741 < NUM_CELL; loop_741++) begin
         if ({b[5],a[23]}) == loop_741[1:0]) begin
          match_flag_741 = 1'b1;
          addr[741] = loop_741[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_742 = 1'b0;
        addr[742] = 3'b0;
        for (loop_742 = 0; loop_742 < NUM_CELL; loop_742++) begin
         if ({b[6],a[23]}) == loop_742[1:0]) begin
          match_flag_742 = 1'b1;
          addr[742] = loop_742[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_743 = 1'b0;
        addr[743] = 3'b0;
        for (loop_743 = 0; loop_743 < NUM_CELL; loop_743++) begin
         if ({b[7],a[23]}) == loop_743[1:0]) begin
          match_flag_743 = 1'b1;
          addr[743] = loop_743[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_744 = 1'b0;
        addr[744] = 3'b0;
        for (loop_744 = 0; loop_744 < NUM_CELL; loop_744++) begin
         if ({b[8],a[23]}) == loop_744[1:0]) begin
          match_flag_744 = 1'b1;
          addr[744] = loop_744[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_745 = 1'b0;
        addr[745] = 3'b0;
        for (loop_745 = 0; loop_745 < NUM_CELL; loop_745++) begin
         if ({b[9],a[23]}) == loop_745[1:0]) begin
          match_flag_745 = 1'b1;
          addr[745] = loop_745[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_746 = 1'b0;
        addr[746] = 3'b0;
        for (loop_746 = 0; loop_746 < NUM_CELL; loop_746++) begin
         if ({b[10],a[23]}) == loop_746[1:0]) begin
          match_flag_746 = 1'b1;
          addr[746] = loop_746[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_747 = 1'b0;
        addr[747] = 3'b0;
        for (loop_747 = 0; loop_747 < NUM_CELL; loop_747++) begin
         if ({b[11],a[23]}) == loop_747[1:0]) begin
          match_flag_747 = 1'b1;
          addr[747] = loop_747[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_748 = 1'b0;
        addr[748] = 3'b0;
        for (loop_748 = 0; loop_748 < NUM_CELL; loop_748++) begin
         if ({b[12],a[23]}) == loop_748[1:0]) begin
          match_flag_748 = 1'b1;
          addr[748] = loop_748[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_749 = 1'b0;
        addr[749] = 3'b0;
        for (loop_749 = 0; loop_749 < NUM_CELL; loop_749++) begin
         if ({b[13],a[23]}) == loop_749[1:0]) begin
          match_flag_749 = 1'b1;
          addr[749] = loop_749[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_750 = 1'b0;
        addr[750] = 3'b0;
        for (loop_750 = 0; loop_750 < NUM_CELL; loop_750++) begin
         if ({b[14],a[23]}) == loop_750[1:0]) begin
          match_flag_750 = 1'b1;
          addr[750] = loop_750[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_751 = 1'b0;
        addr[751] = 3'b0;
        for (loop_751 = 0; loop_751 < NUM_CELL; loop_751++) begin
         if ({b[15],a[23]}) == loop_751[1:0]) begin
          match_flag_751 = 1'b1;
          addr[751] = loop_751[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_752 = 1'b0;
        addr[752] = 3'b0;
        for (loop_752 = 0; loop_752 < NUM_CELL; loop_752++) begin
         if ({b[16],a[23]}) == loop_752[1:0]) begin
          match_flag_752 = 1'b1;
          addr[752] = loop_752[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_753 = 1'b0;
        addr[753] = 3'b0;
        for (loop_753 = 0; loop_753 < NUM_CELL; loop_753++) begin
         if ({b[17],a[23]}) == loop_753[1:0]) begin
          match_flag_753 = 1'b1;
          addr[753] = loop_753[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_754 = 1'b0;
        addr[754] = 3'b0;
        for (loop_754 = 0; loop_754 < NUM_CELL; loop_754++) begin
         if ({b[18],a[23]}) == loop_754[1:0]) begin
          match_flag_754 = 1'b1;
          addr[754] = loop_754[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_755 = 1'b0;
        addr[755] = 3'b0;
        for (loop_755 = 0; loop_755 < NUM_CELL; loop_755++) begin
         if ({b[19],a[23]}) == loop_755[1:0]) begin
          match_flag_755 = 1'b1;
          addr[755] = loop_755[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_756 = 1'b0;
        addr[756] = 3'b0;
        for (loop_756 = 0; loop_756 < NUM_CELL; loop_756++) begin
         if ({b[20],a[23]}) == loop_756[1:0]) begin
          match_flag_756 = 1'b1;
          addr[756] = loop_756[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_757 = 1'b0;
        addr[757] = 3'b0;
        for (loop_757 = 0; loop_757 < NUM_CELL; loop_757++) begin
         if ({b[21],a[23]}) == loop_757[1:0]) begin
          match_flag_757 = 1'b1;
          addr[757] = loop_757[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_758 = 1'b0;
        addr[758] = 3'b0;
        for (loop_758 = 0; loop_758 < NUM_CELL; loop_758++) begin
         if ({b[22],a[23]}) == loop_758[1:0]) begin
          match_flag_758 = 1'b1;
          addr[758] = loop_758[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_759 = 1'b0;
        addr[759] = 3'b0;
        for (loop_759 = 0; loop_759 < NUM_CELL; loop_759++) begin
         if ({b[23],a[23]}) == loop_759[1:0]) begin
          match_flag_759 = 1'b1;
          addr[759] = loop_759[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_760 = 1'b0;
        addr[760] = 3'b0;
        for (loop_760 = 0; loop_760 < NUM_CELL; loop_760++) begin
         if ({b[24],a[23]}) == loop_760[1:0]) begin
          match_flag_760 = 1'b1;
          addr[760] = loop_760[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_761 = 1'b0;
        addr[761] = 3'b0;
        for (loop_761 = 0; loop_761 < NUM_CELL; loop_761++) begin
         if ({b[25],a[23]}) == loop_761[1:0]) begin
          match_flag_761 = 1'b1;
          addr[761] = loop_761[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_762 = 1'b0;
        addr[762] = 3'b0;
        for (loop_762 = 0; loop_762 < NUM_CELL; loop_762++) begin
         if ({b[26],a[23]}) == loop_762[1:0]) begin
          match_flag_762 = 1'b1;
          addr[762] = loop_762[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_763 = 1'b0;
        addr[763] = 3'b0;
        for (loop_763 = 0; loop_763 < NUM_CELL; loop_763++) begin
         if ({b[27],a[23]}) == loop_763[1:0]) begin
          match_flag_763 = 1'b1;
          addr[763] = loop_763[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_764 = 1'b0;
        addr[764] = 3'b0;
        for (loop_764 = 0; loop_764 < NUM_CELL; loop_764++) begin
         if ({b[28],a[23]}) == loop_764[1:0]) begin
          match_flag_764 = 1'b1;
          addr[764] = loop_764[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_765 = 1'b0;
        addr[765] = 3'b0;
        for (loop_765 = 0; loop_765 < NUM_CELL; loop_765++) begin
         if ({b[29],a[23]}) == loop_765[1:0]) begin
          match_flag_765 = 1'b1;
          addr[765] = loop_765[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_766 = 1'b0;
        addr[766] = 3'b0;
        for (loop_766 = 0; loop_766 < NUM_CELL; loop_766++) begin
         if ({b[30],a[23]}) == loop_766[1:0]) begin
          match_flag_766 = 1'b1;
          addr[766] = loop_766[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_767 = 1'b0;
        addr[767] = 3'b0;
        for (loop_767 = 0; loop_767 < NUM_CELL; loop_767++) begin
         if ({b[31],a[23]}) == loop_767[1:0]) begin
          match_flag_767 = 1'b1;
          addr[767] = loop_767[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_768 = 1'b0;
        addr[768] = 3'b0;
        for (loop_768 = 0; loop_768 < NUM_CELL; loop_768++) begin
         if ({b[0],a[24]}) == loop_768[1:0]) begin
          match_flag_768 = 1'b1;
          addr[768] = loop_768[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_769 = 1'b0;
        addr[769] = 3'b0;
        for (loop_769 = 0; loop_769 < NUM_CELL; loop_769++) begin
         if ({b[1],a[24]}) == loop_769[1:0]) begin
          match_flag_769 = 1'b1;
          addr[769] = loop_769[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_770 = 1'b0;
        addr[770] = 3'b0;
        for (loop_770 = 0; loop_770 < NUM_CELL; loop_770++) begin
         if ({b[2],a[24]}) == loop_770[1:0]) begin
          match_flag_770 = 1'b1;
          addr[770] = loop_770[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_771 = 1'b0;
        addr[771] = 3'b0;
        for (loop_771 = 0; loop_771 < NUM_CELL; loop_771++) begin
         if ({b[3],a[24]}) == loop_771[1:0]) begin
          match_flag_771 = 1'b1;
          addr[771] = loop_771[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_772 = 1'b0;
        addr[772] = 3'b0;
        for (loop_772 = 0; loop_772 < NUM_CELL; loop_772++) begin
         if ({b[4],a[24]}) == loop_772[1:0]) begin
          match_flag_772 = 1'b1;
          addr[772] = loop_772[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_773 = 1'b0;
        addr[773] = 3'b0;
        for (loop_773 = 0; loop_773 < NUM_CELL; loop_773++) begin
         if ({b[5],a[24]}) == loop_773[1:0]) begin
          match_flag_773 = 1'b1;
          addr[773] = loop_773[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_774 = 1'b0;
        addr[774] = 3'b0;
        for (loop_774 = 0; loop_774 < NUM_CELL; loop_774++) begin
         if ({b[6],a[24]}) == loop_774[1:0]) begin
          match_flag_774 = 1'b1;
          addr[774] = loop_774[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_775 = 1'b0;
        addr[775] = 3'b0;
        for (loop_775 = 0; loop_775 < NUM_CELL; loop_775++) begin
         if ({b[7],a[24]}) == loop_775[1:0]) begin
          match_flag_775 = 1'b1;
          addr[775] = loop_775[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_776 = 1'b0;
        addr[776] = 3'b0;
        for (loop_776 = 0; loop_776 < NUM_CELL; loop_776++) begin
         if ({b[8],a[24]}) == loop_776[1:0]) begin
          match_flag_776 = 1'b1;
          addr[776] = loop_776[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_777 = 1'b0;
        addr[777] = 3'b0;
        for (loop_777 = 0; loop_777 < NUM_CELL; loop_777++) begin
         if ({b[9],a[24]}) == loop_777[1:0]) begin
          match_flag_777 = 1'b1;
          addr[777] = loop_777[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_778 = 1'b0;
        addr[778] = 3'b0;
        for (loop_778 = 0; loop_778 < NUM_CELL; loop_778++) begin
         if ({b[10],a[24]}) == loop_778[1:0]) begin
          match_flag_778 = 1'b1;
          addr[778] = loop_778[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_779 = 1'b0;
        addr[779] = 3'b0;
        for (loop_779 = 0; loop_779 < NUM_CELL; loop_779++) begin
         if ({b[11],a[24]}) == loop_779[1:0]) begin
          match_flag_779 = 1'b1;
          addr[779] = loop_779[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_780 = 1'b0;
        addr[780] = 3'b0;
        for (loop_780 = 0; loop_780 < NUM_CELL; loop_780++) begin
         if ({b[12],a[24]}) == loop_780[1:0]) begin
          match_flag_780 = 1'b1;
          addr[780] = loop_780[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_781 = 1'b0;
        addr[781] = 3'b0;
        for (loop_781 = 0; loop_781 < NUM_CELL; loop_781++) begin
         if ({b[13],a[24]}) == loop_781[1:0]) begin
          match_flag_781 = 1'b1;
          addr[781] = loop_781[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_782 = 1'b0;
        addr[782] = 3'b0;
        for (loop_782 = 0; loop_782 < NUM_CELL; loop_782++) begin
         if ({b[14],a[24]}) == loop_782[1:0]) begin
          match_flag_782 = 1'b1;
          addr[782] = loop_782[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_783 = 1'b0;
        addr[783] = 3'b0;
        for (loop_783 = 0; loop_783 < NUM_CELL; loop_783++) begin
         if ({b[15],a[24]}) == loop_783[1:0]) begin
          match_flag_783 = 1'b1;
          addr[783] = loop_783[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_784 = 1'b0;
        addr[784] = 3'b0;
        for (loop_784 = 0; loop_784 < NUM_CELL; loop_784++) begin
         if ({b[16],a[24]}) == loop_784[1:0]) begin
          match_flag_784 = 1'b1;
          addr[784] = loop_784[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_785 = 1'b0;
        addr[785] = 3'b0;
        for (loop_785 = 0; loop_785 < NUM_CELL; loop_785++) begin
         if ({b[17],a[24]}) == loop_785[1:0]) begin
          match_flag_785 = 1'b1;
          addr[785] = loop_785[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_786 = 1'b0;
        addr[786] = 3'b0;
        for (loop_786 = 0; loop_786 < NUM_CELL; loop_786++) begin
         if ({b[18],a[24]}) == loop_786[1:0]) begin
          match_flag_786 = 1'b1;
          addr[786] = loop_786[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_787 = 1'b0;
        addr[787] = 3'b0;
        for (loop_787 = 0; loop_787 < NUM_CELL; loop_787++) begin
         if ({b[19],a[24]}) == loop_787[1:0]) begin
          match_flag_787 = 1'b1;
          addr[787] = loop_787[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_788 = 1'b0;
        addr[788] = 3'b0;
        for (loop_788 = 0; loop_788 < NUM_CELL; loop_788++) begin
         if ({b[20],a[24]}) == loop_788[1:0]) begin
          match_flag_788 = 1'b1;
          addr[788] = loop_788[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_789 = 1'b0;
        addr[789] = 3'b0;
        for (loop_789 = 0; loop_789 < NUM_CELL; loop_789++) begin
         if ({b[21],a[24]}) == loop_789[1:0]) begin
          match_flag_789 = 1'b1;
          addr[789] = loop_789[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_790 = 1'b0;
        addr[790] = 3'b0;
        for (loop_790 = 0; loop_790 < NUM_CELL; loop_790++) begin
         if ({b[22],a[24]}) == loop_790[1:0]) begin
          match_flag_790 = 1'b1;
          addr[790] = loop_790[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_791 = 1'b0;
        addr[791] = 3'b0;
        for (loop_791 = 0; loop_791 < NUM_CELL; loop_791++) begin
         if ({b[23],a[24]}) == loop_791[1:0]) begin
          match_flag_791 = 1'b1;
          addr[791] = loop_791[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_792 = 1'b0;
        addr[792] = 3'b0;
        for (loop_792 = 0; loop_792 < NUM_CELL; loop_792++) begin
         if ({b[24],a[24]}) == loop_792[1:0]) begin
          match_flag_792 = 1'b1;
          addr[792] = loop_792[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_793 = 1'b0;
        addr[793] = 3'b0;
        for (loop_793 = 0; loop_793 < NUM_CELL; loop_793++) begin
         if ({b[25],a[24]}) == loop_793[1:0]) begin
          match_flag_793 = 1'b1;
          addr[793] = loop_793[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_794 = 1'b0;
        addr[794] = 3'b0;
        for (loop_794 = 0; loop_794 < NUM_CELL; loop_794++) begin
         if ({b[26],a[24]}) == loop_794[1:0]) begin
          match_flag_794 = 1'b1;
          addr[794] = loop_794[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_795 = 1'b0;
        addr[795] = 3'b0;
        for (loop_795 = 0; loop_795 < NUM_CELL; loop_795++) begin
         if ({b[27],a[24]}) == loop_795[1:0]) begin
          match_flag_795 = 1'b1;
          addr[795] = loop_795[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_796 = 1'b0;
        addr[796] = 3'b0;
        for (loop_796 = 0; loop_796 < NUM_CELL; loop_796++) begin
         if ({b[28],a[24]}) == loop_796[1:0]) begin
          match_flag_796 = 1'b1;
          addr[796] = loop_796[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_797 = 1'b0;
        addr[797] = 3'b0;
        for (loop_797 = 0; loop_797 < NUM_CELL; loop_797++) begin
         if ({b[29],a[24]}) == loop_797[1:0]) begin
          match_flag_797 = 1'b1;
          addr[797] = loop_797[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_798 = 1'b0;
        addr[798] = 3'b0;
        for (loop_798 = 0; loop_798 < NUM_CELL; loop_798++) begin
         if ({b[30],a[24]}) == loop_798[1:0]) begin
          match_flag_798 = 1'b1;
          addr[798] = loop_798[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_799 = 1'b0;
        addr[799] = 3'b0;
        for (loop_799 = 0; loop_799 < NUM_CELL; loop_799++) begin
         if ({b[31],a[24]}) == loop_799[1:0]) begin
          match_flag_799 = 1'b1;
          addr[799] = loop_799[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_800 = 1'b0;
        addr[800] = 3'b0;
        for (loop_800 = 0; loop_800 < NUM_CELL; loop_800++) begin
         if ({b[0],a[25]}) == loop_800[1:0]) begin
          match_flag_800 = 1'b1;
          addr[800] = loop_800[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_801 = 1'b0;
        addr[801] = 3'b0;
        for (loop_801 = 0; loop_801 < NUM_CELL; loop_801++) begin
         if ({b[1],a[25]}) == loop_801[1:0]) begin
          match_flag_801 = 1'b1;
          addr[801] = loop_801[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_802 = 1'b0;
        addr[802] = 3'b0;
        for (loop_802 = 0; loop_802 < NUM_CELL; loop_802++) begin
         if ({b[2],a[25]}) == loop_802[1:0]) begin
          match_flag_802 = 1'b1;
          addr[802] = loop_802[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_803 = 1'b0;
        addr[803] = 3'b0;
        for (loop_803 = 0; loop_803 < NUM_CELL; loop_803++) begin
         if ({b[3],a[25]}) == loop_803[1:0]) begin
          match_flag_803 = 1'b1;
          addr[803] = loop_803[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_804 = 1'b0;
        addr[804] = 3'b0;
        for (loop_804 = 0; loop_804 < NUM_CELL; loop_804++) begin
         if ({b[4],a[25]}) == loop_804[1:0]) begin
          match_flag_804 = 1'b1;
          addr[804] = loop_804[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_805 = 1'b0;
        addr[805] = 3'b0;
        for (loop_805 = 0; loop_805 < NUM_CELL; loop_805++) begin
         if ({b[5],a[25]}) == loop_805[1:0]) begin
          match_flag_805 = 1'b1;
          addr[805] = loop_805[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_806 = 1'b0;
        addr[806] = 3'b0;
        for (loop_806 = 0; loop_806 < NUM_CELL; loop_806++) begin
         if ({b[6],a[25]}) == loop_806[1:0]) begin
          match_flag_806 = 1'b1;
          addr[806] = loop_806[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_807 = 1'b0;
        addr[807] = 3'b0;
        for (loop_807 = 0; loop_807 < NUM_CELL; loop_807++) begin
         if ({b[7],a[25]}) == loop_807[1:0]) begin
          match_flag_807 = 1'b1;
          addr[807] = loop_807[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_808 = 1'b0;
        addr[808] = 3'b0;
        for (loop_808 = 0; loop_808 < NUM_CELL; loop_808++) begin
         if ({b[8],a[25]}) == loop_808[1:0]) begin
          match_flag_808 = 1'b1;
          addr[808] = loop_808[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_809 = 1'b0;
        addr[809] = 3'b0;
        for (loop_809 = 0; loop_809 < NUM_CELL; loop_809++) begin
         if ({b[9],a[25]}) == loop_809[1:0]) begin
          match_flag_809 = 1'b1;
          addr[809] = loop_809[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_810 = 1'b0;
        addr[810] = 3'b0;
        for (loop_810 = 0; loop_810 < NUM_CELL; loop_810++) begin
         if ({b[10],a[25]}) == loop_810[1:0]) begin
          match_flag_810 = 1'b1;
          addr[810] = loop_810[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_811 = 1'b0;
        addr[811] = 3'b0;
        for (loop_811 = 0; loop_811 < NUM_CELL; loop_811++) begin
         if ({b[11],a[25]}) == loop_811[1:0]) begin
          match_flag_811 = 1'b1;
          addr[811] = loop_811[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_812 = 1'b0;
        addr[812] = 3'b0;
        for (loop_812 = 0; loop_812 < NUM_CELL; loop_812++) begin
         if ({b[12],a[25]}) == loop_812[1:0]) begin
          match_flag_812 = 1'b1;
          addr[812] = loop_812[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_813 = 1'b0;
        addr[813] = 3'b0;
        for (loop_813 = 0; loop_813 < NUM_CELL; loop_813++) begin
         if ({b[13],a[25]}) == loop_813[1:0]) begin
          match_flag_813 = 1'b1;
          addr[813] = loop_813[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_814 = 1'b0;
        addr[814] = 3'b0;
        for (loop_814 = 0; loop_814 < NUM_CELL; loop_814++) begin
         if ({b[14],a[25]}) == loop_814[1:0]) begin
          match_flag_814 = 1'b1;
          addr[814] = loop_814[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_815 = 1'b0;
        addr[815] = 3'b0;
        for (loop_815 = 0; loop_815 < NUM_CELL; loop_815++) begin
         if ({b[15],a[25]}) == loop_815[1:0]) begin
          match_flag_815 = 1'b1;
          addr[815] = loop_815[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_816 = 1'b0;
        addr[816] = 3'b0;
        for (loop_816 = 0; loop_816 < NUM_CELL; loop_816++) begin
         if ({b[16],a[25]}) == loop_816[1:0]) begin
          match_flag_816 = 1'b1;
          addr[816] = loop_816[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_817 = 1'b0;
        addr[817] = 3'b0;
        for (loop_817 = 0; loop_817 < NUM_CELL; loop_817++) begin
         if ({b[17],a[25]}) == loop_817[1:0]) begin
          match_flag_817 = 1'b1;
          addr[817] = loop_817[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_818 = 1'b0;
        addr[818] = 3'b0;
        for (loop_818 = 0; loop_818 < NUM_CELL; loop_818++) begin
         if ({b[18],a[25]}) == loop_818[1:0]) begin
          match_flag_818 = 1'b1;
          addr[818] = loop_818[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_819 = 1'b0;
        addr[819] = 3'b0;
        for (loop_819 = 0; loop_819 < NUM_CELL; loop_819++) begin
         if ({b[19],a[25]}) == loop_819[1:0]) begin
          match_flag_819 = 1'b1;
          addr[819] = loop_819[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_820 = 1'b0;
        addr[820] = 3'b0;
        for (loop_820 = 0; loop_820 < NUM_CELL; loop_820++) begin
         if ({b[20],a[25]}) == loop_820[1:0]) begin
          match_flag_820 = 1'b1;
          addr[820] = loop_820[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_821 = 1'b0;
        addr[821] = 3'b0;
        for (loop_821 = 0; loop_821 < NUM_CELL; loop_821++) begin
         if ({b[21],a[25]}) == loop_821[1:0]) begin
          match_flag_821 = 1'b1;
          addr[821] = loop_821[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_822 = 1'b0;
        addr[822] = 3'b0;
        for (loop_822 = 0; loop_822 < NUM_CELL; loop_822++) begin
         if ({b[22],a[25]}) == loop_822[1:0]) begin
          match_flag_822 = 1'b1;
          addr[822] = loop_822[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_823 = 1'b0;
        addr[823] = 3'b0;
        for (loop_823 = 0; loop_823 < NUM_CELL; loop_823++) begin
         if ({b[23],a[25]}) == loop_823[1:0]) begin
          match_flag_823 = 1'b1;
          addr[823] = loop_823[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_824 = 1'b0;
        addr[824] = 3'b0;
        for (loop_824 = 0; loop_824 < NUM_CELL; loop_824++) begin
         if ({b[24],a[25]}) == loop_824[1:0]) begin
          match_flag_824 = 1'b1;
          addr[824] = loop_824[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_825 = 1'b0;
        addr[825] = 3'b0;
        for (loop_825 = 0; loop_825 < NUM_CELL; loop_825++) begin
         if ({b[25],a[25]}) == loop_825[1:0]) begin
          match_flag_825 = 1'b1;
          addr[825] = loop_825[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_826 = 1'b0;
        addr[826] = 3'b0;
        for (loop_826 = 0; loop_826 < NUM_CELL; loop_826++) begin
         if ({b[26],a[25]}) == loop_826[1:0]) begin
          match_flag_826 = 1'b1;
          addr[826] = loop_826[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_827 = 1'b0;
        addr[827] = 3'b0;
        for (loop_827 = 0; loop_827 < NUM_CELL; loop_827++) begin
         if ({b[27],a[25]}) == loop_827[1:0]) begin
          match_flag_827 = 1'b1;
          addr[827] = loop_827[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_828 = 1'b0;
        addr[828] = 3'b0;
        for (loop_828 = 0; loop_828 < NUM_CELL; loop_828++) begin
         if ({b[28],a[25]}) == loop_828[1:0]) begin
          match_flag_828 = 1'b1;
          addr[828] = loop_828[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_829 = 1'b0;
        addr[829] = 3'b0;
        for (loop_829 = 0; loop_829 < NUM_CELL; loop_829++) begin
         if ({b[29],a[25]}) == loop_829[1:0]) begin
          match_flag_829 = 1'b1;
          addr[829] = loop_829[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_830 = 1'b0;
        addr[830] = 3'b0;
        for (loop_830 = 0; loop_830 < NUM_CELL; loop_830++) begin
         if ({b[30],a[25]}) == loop_830[1:0]) begin
          match_flag_830 = 1'b1;
          addr[830] = loop_830[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_831 = 1'b0;
        addr[831] = 3'b0;
        for (loop_831 = 0; loop_831 < NUM_CELL; loop_831++) begin
         if ({b[31],a[25]}) == loop_831[1:0]) begin
          match_flag_831 = 1'b1;
          addr[831] = loop_831[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_832 = 1'b0;
        addr[832] = 3'b0;
        for (loop_832 = 0; loop_832 < NUM_CELL; loop_832++) begin
         if ({b[0],a[26]}) == loop_832[1:0]) begin
          match_flag_832 = 1'b1;
          addr[832] = loop_832[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_833 = 1'b0;
        addr[833] = 3'b0;
        for (loop_833 = 0; loop_833 < NUM_CELL; loop_833++) begin
         if ({b[1],a[26]}) == loop_833[1:0]) begin
          match_flag_833 = 1'b1;
          addr[833] = loop_833[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_834 = 1'b0;
        addr[834] = 3'b0;
        for (loop_834 = 0; loop_834 < NUM_CELL; loop_834++) begin
         if ({b[2],a[26]}) == loop_834[1:0]) begin
          match_flag_834 = 1'b1;
          addr[834] = loop_834[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_835 = 1'b0;
        addr[835] = 3'b0;
        for (loop_835 = 0; loop_835 < NUM_CELL; loop_835++) begin
         if ({b[3],a[26]}) == loop_835[1:0]) begin
          match_flag_835 = 1'b1;
          addr[835] = loop_835[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_836 = 1'b0;
        addr[836] = 3'b0;
        for (loop_836 = 0; loop_836 < NUM_CELL; loop_836++) begin
         if ({b[4],a[26]}) == loop_836[1:0]) begin
          match_flag_836 = 1'b1;
          addr[836] = loop_836[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_837 = 1'b0;
        addr[837] = 3'b0;
        for (loop_837 = 0; loop_837 < NUM_CELL; loop_837++) begin
         if ({b[5],a[26]}) == loop_837[1:0]) begin
          match_flag_837 = 1'b1;
          addr[837] = loop_837[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_838 = 1'b0;
        addr[838] = 3'b0;
        for (loop_838 = 0; loop_838 < NUM_CELL; loop_838++) begin
         if ({b[6],a[26]}) == loop_838[1:0]) begin
          match_flag_838 = 1'b1;
          addr[838] = loop_838[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_839 = 1'b0;
        addr[839] = 3'b0;
        for (loop_839 = 0; loop_839 < NUM_CELL; loop_839++) begin
         if ({b[7],a[26]}) == loop_839[1:0]) begin
          match_flag_839 = 1'b1;
          addr[839] = loop_839[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_840 = 1'b0;
        addr[840] = 3'b0;
        for (loop_840 = 0; loop_840 < NUM_CELL; loop_840++) begin
         if ({b[8],a[26]}) == loop_840[1:0]) begin
          match_flag_840 = 1'b1;
          addr[840] = loop_840[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_841 = 1'b0;
        addr[841] = 3'b0;
        for (loop_841 = 0; loop_841 < NUM_CELL; loop_841++) begin
         if ({b[9],a[26]}) == loop_841[1:0]) begin
          match_flag_841 = 1'b1;
          addr[841] = loop_841[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_842 = 1'b0;
        addr[842] = 3'b0;
        for (loop_842 = 0; loop_842 < NUM_CELL; loop_842++) begin
         if ({b[10],a[26]}) == loop_842[1:0]) begin
          match_flag_842 = 1'b1;
          addr[842] = loop_842[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_843 = 1'b0;
        addr[843] = 3'b0;
        for (loop_843 = 0; loop_843 < NUM_CELL; loop_843++) begin
         if ({b[11],a[26]}) == loop_843[1:0]) begin
          match_flag_843 = 1'b1;
          addr[843] = loop_843[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_844 = 1'b0;
        addr[844] = 3'b0;
        for (loop_844 = 0; loop_844 < NUM_CELL; loop_844++) begin
         if ({b[12],a[26]}) == loop_844[1:0]) begin
          match_flag_844 = 1'b1;
          addr[844] = loop_844[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_845 = 1'b0;
        addr[845] = 3'b0;
        for (loop_845 = 0; loop_845 < NUM_CELL; loop_845++) begin
         if ({b[13],a[26]}) == loop_845[1:0]) begin
          match_flag_845 = 1'b1;
          addr[845] = loop_845[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_846 = 1'b0;
        addr[846] = 3'b0;
        for (loop_846 = 0; loop_846 < NUM_CELL; loop_846++) begin
         if ({b[14],a[26]}) == loop_846[1:0]) begin
          match_flag_846 = 1'b1;
          addr[846] = loop_846[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_847 = 1'b0;
        addr[847] = 3'b0;
        for (loop_847 = 0; loop_847 < NUM_CELL; loop_847++) begin
         if ({b[15],a[26]}) == loop_847[1:0]) begin
          match_flag_847 = 1'b1;
          addr[847] = loop_847[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_848 = 1'b0;
        addr[848] = 3'b0;
        for (loop_848 = 0; loop_848 < NUM_CELL; loop_848++) begin
         if ({b[16],a[26]}) == loop_848[1:0]) begin
          match_flag_848 = 1'b1;
          addr[848] = loop_848[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_849 = 1'b0;
        addr[849] = 3'b0;
        for (loop_849 = 0; loop_849 < NUM_CELL; loop_849++) begin
         if ({b[17],a[26]}) == loop_849[1:0]) begin
          match_flag_849 = 1'b1;
          addr[849] = loop_849[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_850 = 1'b0;
        addr[850] = 3'b0;
        for (loop_850 = 0; loop_850 < NUM_CELL; loop_850++) begin
         if ({b[18],a[26]}) == loop_850[1:0]) begin
          match_flag_850 = 1'b1;
          addr[850] = loop_850[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_851 = 1'b0;
        addr[851] = 3'b0;
        for (loop_851 = 0; loop_851 < NUM_CELL; loop_851++) begin
         if ({b[19],a[26]}) == loop_851[1:0]) begin
          match_flag_851 = 1'b1;
          addr[851] = loop_851[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_852 = 1'b0;
        addr[852] = 3'b0;
        for (loop_852 = 0; loop_852 < NUM_CELL; loop_852++) begin
         if ({b[20],a[26]}) == loop_852[1:0]) begin
          match_flag_852 = 1'b1;
          addr[852] = loop_852[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_853 = 1'b0;
        addr[853] = 3'b0;
        for (loop_853 = 0; loop_853 < NUM_CELL; loop_853++) begin
         if ({b[21],a[26]}) == loop_853[1:0]) begin
          match_flag_853 = 1'b1;
          addr[853] = loop_853[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_854 = 1'b0;
        addr[854] = 3'b0;
        for (loop_854 = 0; loop_854 < NUM_CELL; loop_854++) begin
         if ({b[22],a[26]}) == loop_854[1:0]) begin
          match_flag_854 = 1'b1;
          addr[854] = loop_854[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_855 = 1'b0;
        addr[855] = 3'b0;
        for (loop_855 = 0; loop_855 < NUM_CELL; loop_855++) begin
         if ({b[23],a[26]}) == loop_855[1:0]) begin
          match_flag_855 = 1'b1;
          addr[855] = loop_855[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_856 = 1'b0;
        addr[856] = 3'b0;
        for (loop_856 = 0; loop_856 < NUM_CELL; loop_856++) begin
         if ({b[24],a[26]}) == loop_856[1:0]) begin
          match_flag_856 = 1'b1;
          addr[856] = loop_856[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_857 = 1'b0;
        addr[857] = 3'b0;
        for (loop_857 = 0; loop_857 < NUM_CELL; loop_857++) begin
         if ({b[25],a[26]}) == loop_857[1:0]) begin
          match_flag_857 = 1'b1;
          addr[857] = loop_857[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_858 = 1'b0;
        addr[858] = 3'b0;
        for (loop_858 = 0; loop_858 < NUM_CELL; loop_858++) begin
         if ({b[26],a[26]}) == loop_858[1:0]) begin
          match_flag_858 = 1'b1;
          addr[858] = loop_858[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_859 = 1'b0;
        addr[859] = 3'b0;
        for (loop_859 = 0; loop_859 < NUM_CELL; loop_859++) begin
         if ({b[27],a[26]}) == loop_859[1:0]) begin
          match_flag_859 = 1'b1;
          addr[859] = loop_859[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_860 = 1'b0;
        addr[860] = 3'b0;
        for (loop_860 = 0; loop_860 < NUM_CELL; loop_860++) begin
         if ({b[28],a[26]}) == loop_860[1:0]) begin
          match_flag_860 = 1'b1;
          addr[860] = loop_860[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_861 = 1'b0;
        addr[861] = 3'b0;
        for (loop_861 = 0; loop_861 < NUM_CELL; loop_861++) begin
         if ({b[29],a[26]}) == loop_861[1:0]) begin
          match_flag_861 = 1'b1;
          addr[861] = loop_861[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_862 = 1'b0;
        addr[862] = 3'b0;
        for (loop_862 = 0; loop_862 < NUM_CELL; loop_862++) begin
         if ({b[30],a[26]}) == loop_862[1:0]) begin
          match_flag_862 = 1'b1;
          addr[862] = loop_862[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_863 = 1'b0;
        addr[863] = 3'b0;
        for (loop_863 = 0; loop_863 < NUM_CELL; loop_863++) begin
         if ({b[31],a[26]}) == loop_863[1:0]) begin
          match_flag_863 = 1'b1;
          addr[863] = loop_863[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_864 = 1'b0;
        addr[864] = 3'b0;
        for (loop_864 = 0; loop_864 < NUM_CELL; loop_864++) begin
         if ({b[0],a[27]}) == loop_864[1:0]) begin
          match_flag_864 = 1'b1;
          addr[864] = loop_864[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_865 = 1'b0;
        addr[865] = 3'b0;
        for (loop_865 = 0; loop_865 < NUM_CELL; loop_865++) begin
         if ({b[1],a[27]}) == loop_865[1:0]) begin
          match_flag_865 = 1'b1;
          addr[865] = loop_865[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_866 = 1'b0;
        addr[866] = 3'b0;
        for (loop_866 = 0; loop_866 < NUM_CELL; loop_866++) begin
         if ({b[2],a[27]}) == loop_866[1:0]) begin
          match_flag_866 = 1'b1;
          addr[866] = loop_866[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_867 = 1'b0;
        addr[867] = 3'b0;
        for (loop_867 = 0; loop_867 < NUM_CELL; loop_867++) begin
         if ({b[3],a[27]}) == loop_867[1:0]) begin
          match_flag_867 = 1'b1;
          addr[867] = loop_867[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_868 = 1'b0;
        addr[868] = 3'b0;
        for (loop_868 = 0; loop_868 < NUM_CELL; loop_868++) begin
         if ({b[4],a[27]}) == loop_868[1:0]) begin
          match_flag_868 = 1'b1;
          addr[868] = loop_868[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_869 = 1'b0;
        addr[869] = 3'b0;
        for (loop_869 = 0; loop_869 < NUM_CELL; loop_869++) begin
         if ({b[5],a[27]}) == loop_869[1:0]) begin
          match_flag_869 = 1'b1;
          addr[869] = loop_869[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_870 = 1'b0;
        addr[870] = 3'b0;
        for (loop_870 = 0; loop_870 < NUM_CELL; loop_870++) begin
         if ({b[6],a[27]}) == loop_870[1:0]) begin
          match_flag_870 = 1'b1;
          addr[870] = loop_870[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_871 = 1'b0;
        addr[871] = 3'b0;
        for (loop_871 = 0; loop_871 < NUM_CELL; loop_871++) begin
         if ({b[7],a[27]}) == loop_871[1:0]) begin
          match_flag_871 = 1'b1;
          addr[871] = loop_871[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_872 = 1'b0;
        addr[872] = 3'b0;
        for (loop_872 = 0; loop_872 < NUM_CELL; loop_872++) begin
         if ({b[8],a[27]}) == loop_872[1:0]) begin
          match_flag_872 = 1'b1;
          addr[872] = loop_872[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_873 = 1'b0;
        addr[873] = 3'b0;
        for (loop_873 = 0; loop_873 < NUM_CELL; loop_873++) begin
         if ({b[9],a[27]}) == loop_873[1:0]) begin
          match_flag_873 = 1'b1;
          addr[873] = loop_873[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_874 = 1'b0;
        addr[874] = 3'b0;
        for (loop_874 = 0; loop_874 < NUM_CELL; loop_874++) begin
         if ({b[10],a[27]}) == loop_874[1:0]) begin
          match_flag_874 = 1'b1;
          addr[874] = loop_874[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_875 = 1'b0;
        addr[875] = 3'b0;
        for (loop_875 = 0; loop_875 < NUM_CELL; loop_875++) begin
         if ({b[11],a[27]}) == loop_875[1:0]) begin
          match_flag_875 = 1'b1;
          addr[875] = loop_875[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_876 = 1'b0;
        addr[876] = 3'b0;
        for (loop_876 = 0; loop_876 < NUM_CELL; loop_876++) begin
         if ({b[12],a[27]}) == loop_876[1:0]) begin
          match_flag_876 = 1'b1;
          addr[876] = loop_876[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_877 = 1'b0;
        addr[877] = 3'b0;
        for (loop_877 = 0; loop_877 < NUM_CELL; loop_877++) begin
         if ({b[13],a[27]}) == loop_877[1:0]) begin
          match_flag_877 = 1'b1;
          addr[877] = loop_877[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_878 = 1'b0;
        addr[878] = 3'b0;
        for (loop_878 = 0; loop_878 < NUM_CELL; loop_878++) begin
         if ({b[14],a[27]}) == loop_878[1:0]) begin
          match_flag_878 = 1'b1;
          addr[878] = loop_878[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_879 = 1'b0;
        addr[879] = 3'b0;
        for (loop_879 = 0; loop_879 < NUM_CELL; loop_879++) begin
         if ({b[15],a[27]}) == loop_879[1:0]) begin
          match_flag_879 = 1'b1;
          addr[879] = loop_879[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_880 = 1'b0;
        addr[880] = 3'b0;
        for (loop_880 = 0; loop_880 < NUM_CELL; loop_880++) begin
         if ({b[16],a[27]}) == loop_880[1:0]) begin
          match_flag_880 = 1'b1;
          addr[880] = loop_880[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_881 = 1'b0;
        addr[881] = 3'b0;
        for (loop_881 = 0; loop_881 < NUM_CELL; loop_881++) begin
         if ({b[17],a[27]}) == loop_881[1:0]) begin
          match_flag_881 = 1'b1;
          addr[881] = loop_881[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_882 = 1'b0;
        addr[882] = 3'b0;
        for (loop_882 = 0; loop_882 < NUM_CELL; loop_882++) begin
         if ({b[18],a[27]}) == loop_882[1:0]) begin
          match_flag_882 = 1'b1;
          addr[882] = loop_882[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_883 = 1'b0;
        addr[883] = 3'b0;
        for (loop_883 = 0; loop_883 < NUM_CELL; loop_883++) begin
         if ({b[19],a[27]}) == loop_883[1:0]) begin
          match_flag_883 = 1'b1;
          addr[883] = loop_883[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_884 = 1'b0;
        addr[884] = 3'b0;
        for (loop_884 = 0; loop_884 < NUM_CELL; loop_884++) begin
         if ({b[20],a[27]}) == loop_884[1:0]) begin
          match_flag_884 = 1'b1;
          addr[884] = loop_884[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_885 = 1'b0;
        addr[885] = 3'b0;
        for (loop_885 = 0; loop_885 < NUM_CELL; loop_885++) begin
         if ({b[21],a[27]}) == loop_885[1:0]) begin
          match_flag_885 = 1'b1;
          addr[885] = loop_885[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_886 = 1'b0;
        addr[886] = 3'b0;
        for (loop_886 = 0; loop_886 < NUM_CELL; loop_886++) begin
         if ({b[22],a[27]}) == loop_886[1:0]) begin
          match_flag_886 = 1'b1;
          addr[886] = loop_886[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_887 = 1'b0;
        addr[887] = 3'b0;
        for (loop_887 = 0; loop_887 < NUM_CELL; loop_887++) begin
         if ({b[23],a[27]}) == loop_887[1:0]) begin
          match_flag_887 = 1'b1;
          addr[887] = loop_887[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_888 = 1'b0;
        addr[888] = 3'b0;
        for (loop_888 = 0; loop_888 < NUM_CELL; loop_888++) begin
         if ({b[24],a[27]}) == loop_888[1:0]) begin
          match_flag_888 = 1'b1;
          addr[888] = loop_888[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_889 = 1'b0;
        addr[889] = 3'b0;
        for (loop_889 = 0; loop_889 < NUM_CELL; loop_889++) begin
         if ({b[25],a[27]}) == loop_889[1:0]) begin
          match_flag_889 = 1'b1;
          addr[889] = loop_889[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_890 = 1'b0;
        addr[890] = 3'b0;
        for (loop_890 = 0; loop_890 < NUM_CELL; loop_890++) begin
         if ({b[26],a[27]}) == loop_890[1:0]) begin
          match_flag_890 = 1'b1;
          addr[890] = loop_890[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_891 = 1'b0;
        addr[891] = 3'b0;
        for (loop_891 = 0; loop_891 < NUM_CELL; loop_891++) begin
         if ({b[27],a[27]}) == loop_891[1:0]) begin
          match_flag_891 = 1'b1;
          addr[891] = loop_891[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_892 = 1'b0;
        addr[892] = 3'b0;
        for (loop_892 = 0; loop_892 < NUM_CELL; loop_892++) begin
         if ({b[28],a[27]}) == loop_892[1:0]) begin
          match_flag_892 = 1'b1;
          addr[892] = loop_892[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_893 = 1'b0;
        addr[893] = 3'b0;
        for (loop_893 = 0; loop_893 < NUM_CELL; loop_893++) begin
         if ({b[29],a[27]}) == loop_893[1:0]) begin
          match_flag_893 = 1'b1;
          addr[893] = loop_893[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_894 = 1'b0;
        addr[894] = 3'b0;
        for (loop_894 = 0; loop_894 < NUM_CELL; loop_894++) begin
         if ({b[30],a[27]}) == loop_894[1:0]) begin
          match_flag_894 = 1'b1;
          addr[894] = loop_894[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_895 = 1'b0;
        addr[895] = 3'b0;
        for (loop_895 = 0; loop_895 < NUM_CELL; loop_895++) begin
         if ({b[31],a[27]}) == loop_895[1:0]) begin
          match_flag_895 = 1'b1;
          addr[895] = loop_895[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_896 = 1'b0;
        addr[896] = 3'b0;
        for (loop_896 = 0; loop_896 < NUM_CELL; loop_896++) begin
         if ({b[0],a[28]}) == loop_896[1:0]) begin
          match_flag_896 = 1'b1;
          addr[896] = loop_896[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_897 = 1'b0;
        addr[897] = 3'b0;
        for (loop_897 = 0; loop_897 < NUM_CELL; loop_897++) begin
         if ({b[1],a[28]}) == loop_897[1:0]) begin
          match_flag_897 = 1'b1;
          addr[897] = loop_897[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_898 = 1'b0;
        addr[898] = 3'b0;
        for (loop_898 = 0; loop_898 < NUM_CELL; loop_898++) begin
         if ({b[2],a[28]}) == loop_898[1:0]) begin
          match_flag_898 = 1'b1;
          addr[898] = loop_898[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_899 = 1'b0;
        addr[899] = 3'b0;
        for (loop_899 = 0; loop_899 < NUM_CELL; loop_899++) begin
         if ({b[3],a[28]}) == loop_899[1:0]) begin
          match_flag_899 = 1'b1;
          addr[899] = loop_899[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_900 = 1'b0;
        addr[900] = 3'b0;
        for (loop_900 = 0; loop_900 < NUM_CELL; loop_900++) begin
         if ({b[4],a[28]}) == loop_900[1:0]) begin
          match_flag_900 = 1'b1;
          addr[900] = loop_900[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_901 = 1'b0;
        addr[901] = 3'b0;
        for (loop_901 = 0; loop_901 < NUM_CELL; loop_901++) begin
         if ({b[5],a[28]}) == loop_901[1:0]) begin
          match_flag_901 = 1'b1;
          addr[901] = loop_901[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_902 = 1'b0;
        addr[902] = 3'b0;
        for (loop_902 = 0; loop_902 < NUM_CELL; loop_902++) begin
         if ({b[6],a[28]}) == loop_902[1:0]) begin
          match_flag_902 = 1'b1;
          addr[902] = loop_902[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_903 = 1'b0;
        addr[903] = 3'b0;
        for (loop_903 = 0; loop_903 < NUM_CELL; loop_903++) begin
         if ({b[7],a[28]}) == loop_903[1:0]) begin
          match_flag_903 = 1'b1;
          addr[903] = loop_903[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_904 = 1'b0;
        addr[904] = 3'b0;
        for (loop_904 = 0; loop_904 < NUM_CELL; loop_904++) begin
         if ({b[8],a[28]}) == loop_904[1:0]) begin
          match_flag_904 = 1'b1;
          addr[904] = loop_904[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_905 = 1'b0;
        addr[905] = 3'b0;
        for (loop_905 = 0; loop_905 < NUM_CELL; loop_905++) begin
         if ({b[9],a[28]}) == loop_905[1:0]) begin
          match_flag_905 = 1'b1;
          addr[905] = loop_905[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_906 = 1'b0;
        addr[906] = 3'b0;
        for (loop_906 = 0; loop_906 < NUM_CELL; loop_906++) begin
         if ({b[10],a[28]}) == loop_906[1:0]) begin
          match_flag_906 = 1'b1;
          addr[906] = loop_906[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_907 = 1'b0;
        addr[907] = 3'b0;
        for (loop_907 = 0; loop_907 < NUM_CELL; loop_907++) begin
         if ({b[11],a[28]}) == loop_907[1:0]) begin
          match_flag_907 = 1'b1;
          addr[907] = loop_907[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_908 = 1'b0;
        addr[908] = 3'b0;
        for (loop_908 = 0; loop_908 < NUM_CELL; loop_908++) begin
         if ({b[12],a[28]}) == loop_908[1:0]) begin
          match_flag_908 = 1'b1;
          addr[908] = loop_908[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_909 = 1'b0;
        addr[909] = 3'b0;
        for (loop_909 = 0; loop_909 < NUM_CELL; loop_909++) begin
         if ({b[13],a[28]}) == loop_909[1:0]) begin
          match_flag_909 = 1'b1;
          addr[909] = loop_909[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_910 = 1'b0;
        addr[910] = 3'b0;
        for (loop_910 = 0; loop_910 < NUM_CELL; loop_910++) begin
         if ({b[14],a[28]}) == loop_910[1:0]) begin
          match_flag_910 = 1'b1;
          addr[910] = loop_910[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_911 = 1'b0;
        addr[911] = 3'b0;
        for (loop_911 = 0; loop_911 < NUM_CELL; loop_911++) begin
         if ({b[15],a[28]}) == loop_911[1:0]) begin
          match_flag_911 = 1'b1;
          addr[911] = loop_911[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_912 = 1'b0;
        addr[912] = 3'b0;
        for (loop_912 = 0; loop_912 < NUM_CELL; loop_912++) begin
         if ({b[16],a[28]}) == loop_912[1:0]) begin
          match_flag_912 = 1'b1;
          addr[912] = loop_912[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_913 = 1'b0;
        addr[913] = 3'b0;
        for (loop_913 = 0; loop_913 < NUM_CELL; loop_913++) begin
         if ({b[17],a[28]}) == loop_913[1:0]) begin
          match_flag_913 = 1'b1;
          addr[913] = loop_913[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_914 = 1'b0;
        addr[914] = 3'b0;
        for (loop_914 = 0; loop_914 < NUM_CELL; loop_914++) begin
         if ({b[18],a[28]}) == loop_914[1:0]) begin
          match_flag_914 = 1'b1;
          addr[914] = loop_914[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_915 = 1'b0;
        addr[915] = 3'b0;
        for (loop_915 = 0; loop_915 < NUM_CELL; loop_915++) begin
         if ({b[19],a[28]}) == loop_915[1:0]) begin
          match_flag_915 = 1'b1;
          addr[915] = loop_915[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_916 = 1'b0;
        addr[916] = 3'b0;
        for (loop_916 = 0; loop_916 < NUM_CELL; loop_916++) begin
         if ({b[20],a[28]}) == loop_916[1:0]) begin
          match_flag_916 = 1'b1;
          addr[916] = loop_916[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_917 = 1'b0;
        addr[917] = 3'b0;
        for (loop_917 = 0; loop_917 < NUM_CELL; loop_917++) begin
         if ({b[21],a[28]}) == loop_917[1:0]) begin
          match_flag_917 = 1'b1;
          addr[917] = loop_917[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_918 = 1'b0;
        addr[918] = 3'b0;
        for (loop_918 = 0; loop_918 < NUM_CELL; loop_918++) begin
         if ({b[22],a[28]}) == loop_918[1:0]) begin
          match_flag_918 = 1'b1;
          addr[918] = loop_918[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_919 = 1'b0;
        addr[919] = 3'b0;
        for (loop_919 = 0; loop_919 < NUM_CELL; loop_919++) begin
         if ({b[23],a[28]}) == loop_919[1:0]) begin
          match_flag_919 = 1'b1;
          addr[919] = loop_919[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_920 = 1'b0;
        addr[920] = 3'b0;
        for (loop_920 = 0; loop_920 < NUM_CELL; loop_920++) begin
         if ({b[24],a[28]}) == loop_920[1:0]) begin
          match_flag_920 = 1'b1;
          addr[920] = loop_920[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_921 = 1'b0;
        addr[921] = 3'b0;
        for (loop_921 = 0; loop_921 < NUM_CELL; loop_921++) begin
         if ({b[25],a[28]}) == loop_921[1:0]) begin
          match_flag_921 = 1'b1;
          addr[921] = loop_921[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_922 = 1'b0;
        addr[922] = 3'b0;
        for (loop_922 = 0; loop_922 < NUM_CELL; loop_922++) begin
         if ({b[26],a[28]}) == loop_922[1:0]) begin
          match_flag_922 = 1'b1;
          addr[922] = loop_922[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_923 = 1'b0;
        addr[923] = 3'b0;
        for (loop_923 = 0; loop_923 < NUM_CELL; loop_923++) begin
         if ({b[27],a[28]}) == loop_923[1:0]) begin
          match_flag_923 = 1'b1;
          addr[923] = loop_923[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_924 = 1'b0;
        addr[924] = 3'b0;
        for (loop_924 = 0; loop_924 < NUM_CELL; loop_924++) begin
         if ({b[28],a[28]}) == loop_924[1:0]) begin
          match_flag_924 = 1'b1;
          addr[924] = loop_924[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_925 = 1'b0;
        addr[925] = 3'b0;
        for (loop_925 = 0; loop_925 < NUM_CELL; loop_925++) begin
         if ({b[29],a[28]}) == loop_925[1:0]) begin
          match_flag_925 = 1'b1;
          addr[925] = loop_925[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_926 = 1'b0;
        addr[926] = 3'b0;
        for (loop_926 = 0; loop_926 < NUM_CELL; loop_926++) begin
         if ({b[30],a[28]}) == loop_926[1:0]) begin
          match_flag_926 = 1'b1;
          addr[926] = loop_926[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_927 = 1'b0;
        addr[927] = 3'b0;
        for (loop_927 = 0; loop_927 < NUM_CELL; loop_927++) begin
         if ({b[31],a[28]}) == loop_927[1:0]) begin
          match_flag_927 = 1'b1;
          addr[927] = loop_927[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_928 = 1'b0;
        addr[928] = 3'b0;
        for (loop_928 = 0; loop_928 < NUM_CELL; loop_928++) begin
         if ({b[0],a[29]}) == loop_928[1:0]) begin
          match_flag_928 = 1'b1;
          addr[928] = loop_928[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_929 = 1'b0;
        addr[929] = 3'b0;
        for (loop_929 = 0; loop_929 < NUM_CELL; loop_929++) begin
         if ({b[1],a[29]}) == loop_929[1:0]) begin
          match_flag_929 = 1'b1;
          addr[929] = loop_929[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_930 = 1'b0;
        addr[930] = 3'b0;
        for (loop_930 = 0; loop_930 < NUM_CELL; loop_930++) begin
         if ({b[2],a[29]}) == loop_930[1:0]) begin
          match_flag_930 = 1'b1;
          addr[930] = loop_930[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_931 = 1'b0;
        addr[931] = 3'b0;
        for (loop_931 = 0; loop_931 < NUM_CELL; loop_931++) begin
         if ({b[3],a[29]}) == loop_931[1:0]) begin
          match_flag_931 = 1'b1;
          addr[931] = loop_931[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_932 = 1'b0;
        addr[932] = 3'b0;
        for (loop_932 = 0; loop_932 < NUM_CELL; loop_932++) begin
         if ({b[4],a[29]}) == loop_932[1:0]) begin
          match_flag_932 = 1'b1;
          addr[932] = loop_932[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_933 = 1'b0;
        addr[933] = 3'b0;
        for (loop_933 = 0; loop_933 < NUM_CELL; loop_933++) begin
         if ({b[5],a[29]}) == loop_933[1:0]) begin
          match_flag_933 = 1'b1;
          addr[933] = loop_933[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_934 = 1'b0;
        addr[934] = 3'b0;
        for (loop_934 = 0; loop_934 < NUM_CELL; loop_934++) begin
         if ({b[6],a[29]}) == loop_934[1:0]) begin
          match_flag_934 = 1'b1;
          addr[934] = loop_934[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_935 = 1'b0;
        addr[935] = 3'b0;
        for (loop_935 = 0; loop_935 < NUM_CELL; loop_935++) begin
         if ({b[7],a[29]}) == loop_935[1:0]) begin
          match_flag_935 = 1'b1;
          addr[935] = loop_935[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_936 = 1'b0;
        addr[936] = 3'b0;
        for (loop_936 = 0; loop_936 < NUM_CELL; loop_936++) begin
         if ({b[8],a[29]}) == loop_936[1:0]) begin
          match_flag_936 = 1'b1;
          addr[936] = loop_936[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_937 = 1'b0;
        addr[937] = 3'b0;
        for (loop_937 = 0; loop_937 < NUM_CELL; loop_937++) begin
         if ({b[9],a[29]}) == loop_937[1:0]) begin
          match_flag_937 = 1'b1;
          addr[937] = loop_937[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_938 = 1'b0;
        addr[938] = 3'b0;
        for (loop_938 = 0; loop_938 < NUM_CELL; loop_938++) begin
         if ({b[10],a[29]}) == loop_938[1:0]) begin
          match_flag_938 = 1'b1;
          addr[938] = loop_938[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_939 = 1'b0;
        addr[939] = 3'b0;
        for (loop_939 = 0; loop_939 < NUM_CELL; loop_939++) begin
         if ({b[11],a[29]}) == loop_939[1:0]) begin
          match_flag_939 = 1'b1;
          addr[939] = loop_939[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_940 = 1'b0;
        addr[940] = 3'b0;
        for (loop_940 = 0; loop_940 < NUM_CELL; loop_940++) begin
         if ({b[12],a[29]}) == loop_940[1:0]) begin
          match_flag_940 = 1'b1;
          addr[940] = loop_940[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_941 = 1'b0;
        addr[941] = 3'b0;
        for (loop_941 = 0; loop_941 < NUM_CELL; loop_941++) begin
         if ({b[13],a[29]}) == loop_941[1:0]) begin
          match_flag_941 = 1'b1;
          addr[941] = loop_941[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_942 = 1'b0;
        addr[942] = 3'b0;
        for (loop_942 = 0; loop_942 < NUM_CELL; loop_942++) begin
         if ({b[14],a[29]}) == loop_942[1:0]) begin
          match_flag_942 = 1'b1;
          addr[942] = loop_942[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_943 = 1'b0;
        addr[943] = 3'b0;
        for (loop_943 = 0; loop_943 < NUM_CELL; loop_943++) begin
         if ({b[15],a[29]}) == loop_943[1:0]) begin
          match_flag_943 = 1'b1;
          addr[943] = loop_943[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_944 = 1'b0;
        addr[944] = 3'b0;
        for (loop_944 = 0; loop_944 < NUM_CELL; loop_944++) begin
         if ({b[16],a[29]}) == loop_944[1:0]) begin
          match_flag_944 = 1'b1;
          addr[944] = loop_944[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_945 = 1'b0;
        addr[945] = 3'b0;
        for (loop_945 = 0; loop_945 < NUM_CELL; loop_945++) begin
         if ({b[17],a[29]}) == loop_945[1:0]) begin
          match_flag_945 = 1'b1;
          addr[945] = loop_945[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_946 = 1'b0;
        addr[946] = 3'b0;
        for (loop_946 = 0; loop_946 < NUM_CELL; loop_946++) begin
         if ({b[18],a[29]}) == loop_946[1:0]) begin
          match_flag_946 = 1'b1;
          addr[946] = loop_946[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_947 = 1'b0;
        addr[947] = 3'b0;
        for (loop_947 = 0; loop_947 < NUM_CELL; loop_947++) begin
         if ({b[19],a[29]}) == loop_947[1:0]) begin
          match_flag_947 = 1'b1;
          addr[947] = loop_947[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_948 = 1'b0;
        addr[948] = 3'b0;
        for (loop_948 = 0; loop_948 < NUM_CELL; loop_948++) begin
         if ({b[20],a[29]}) == loop_948[1:0]) begin
          match_flag_948 = 1'b1;
          addr[948] = loop_948[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_949 = 1'b0;
        addr[949] = 3'b0;
        for (loop_949 = 0; loop_949 < NUM_CELL; loop_949++) begin
         if ({b[21],a[29]}) == loop_949[1:0]) begin
          match_flag_949 = 1'b1;
          addr[949] = loop_949[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_950 = 1'b0;
        addr[950] = 3'b0;
        for (loop_950 = 0; loop_950 < NUM_CELL; loop_950++) begin
         if ({b[22],a[29]}) == loop_950[1:0]) begin
          match_flag_950 = 1'b1;
          addr[950] = loop_950[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_951 = 1'b0;
        addr[951] = 3'b0;
        for (loop_951 = 0; loop_951 < NUM_CELL; loop_951++) begin
         if ({b[23],a[29]}) == loop_951[1:0]) begin
          match_flag_951 = 1'b1;
          addr[951] = loop_951[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_952 = 1'b0;
        addr[952] = 3'b0;
        for (loop_952 = 0; loop_952 < NUM_CELL; loop_952++) begin
         if ({b[24],a[29]}) == loop_952[1:0]) begin
          match_flag_952 = 1'b1;
          addr[952] = loop_952[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_953 = 1'b0;
        addr[953] = 3'b0;
        for (loop_953 = 0; loop_953 < NUM_CELL; loop_953++) begin
         if ({b[25],a[29]}) == loop_953[1:0]) begin
          match_flag_953 = 1'b1;
          addr[953] = loop_953[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_954 = 1'b0;
        addr[954] = 3'b0;
        for (loop_954 = 0; loop_954 < NUM_CELL; loop_954++) begin
         if ({b[26],a[29]}) == loop_954[1:0]) begin
          match_flag_954 = 1'b1;
          addr[954] = loop_954[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_955 = 1'b0;
        addr[955] = 3'b0;
        for (loop_955 = 0; loop_955 < NUM_CELL; loop_955++) begin
         if ({b[27],a[29]}) == loop_955[1:0]) begin
          match_flag_955 = 1'b1;
          addr[955] = loop_955[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_956 = 1'b0;
        addr[956] = 3'b0;
        for (loop_956 = 0; loop_956 < NUM_CELL; loop_956++) begin
         if ({b[28],a[29]}) == loop_956[1:0]) begin
          match_flag_956 = 1'b1;
          addr[956] = loop_956[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_957 = 1'b0;
        addr[957] = 3'b0;
        for (loop_957 = 0; loop_957 < NUM_CELL; loop_957++) begin
         if ({b[29],a[29]}) == loop_957[1:0]) begin
          match_flag_957 = 1'b1;
          addr[957] = loop_957[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_958 = 1'b0;
        addr[958] = 3'b0;
        for (loop_958 = 0; loop_958 < NUM_CELL; loop_958++) begin
         if ({b[30],a[29]}) == loop_958[1:0]) begin
          match_flag_958 = 1'b1;
          addr[958] = loop_958[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_959 = 1'b0;
        addr[959] = 3'b0;
        for (loop_959 = 0; loop_959 < NUM_CELL; loop_959++) begin
         if ({b[31],a[29]}) == loop_959[1:0]) begin
          match_flag_959 = 1'b1;
          addr[959] = loop_959[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_960 = 1'b0;
        addr[960] = 3'b0;
        for (loop_960 = 0; loop_960 < NUM_CELL; loop_960++) begin
         if ({b[0],a[30]}) == loop_960[1:0]) begin
          match_flag_960 = 1'b1;
          addr[960] = loop_960[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_961 = 1'b0;
        addr[961] = 3'b0;
        for (loop_961 = 0; loop_961 < NUM_CELL; loop_961++) begin
         if ({b[1],a[30]}) == loop_961[1:0]) begin
          match_flag_961 = 1'b1;
          addr[961] = loop_961[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_962 = 1'b0;
        addr[962] = 3'b0;
        for (loop_962 = 0; loop_962 < NUM_CELL; loop_962++) begin
         if ({b[2],a[30]}) == loop_962[1:0]) begin
          match_flag_962 = 1'b1;
          addr[962] = loop_962[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_963 = 1'b0;
        addr[963] = 3'b0;
        for (loop_963 = 0; loop_963 < NUM_CELL; loop_963++) begin
         if ({b[3],a[30]}) == loop_963[1:0]) begin
          match_flag_963 = 1'b1;
          addr[963] = loop_963[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_964 = 1'b0;
        addr[964] = 3'b0;
        for (loop_964 = 0; loop_964 < NUM_CELL; loop_964++) begin
         if ({b[4],a[30]}) == loop_964[1:0]) begin
          match_flag_964 = 1'b1;
          addr[964] = loop_964[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_965 = 1'b0;
        addr[965] = 3'b0;
        for (loop_965 = 0; loop_965 < NUM_CELL; loop_965++) begin
         if ({b[5],a[30]}) == loop_965[1:0]) begin
          match_flag_965 = 1'b1;
          addr[965] = loop_965[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_966 = 1'b0;
        addr[966] = 3'b0;
        for (loop_966 = 0; loop_966 < NUM_CELL; loop_966++) begin
         if ({b[6],a[30]}) == loop_966[1:0]) begin
          match_flag_966 = 1'b1;
          addr[966] = loop_966[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_967 = 1'b0;
        addr[967] = 3'b0;
        for (loop_967 = 0; loop_967 < NUM_CELL; loop_967++) begin
         if ({b[7],a[30]}) == loop_967[1:0]) begin
          match_flag_967 = 1'b1;
          addr[967] = loop_967[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_968 = 1'b0;
        addr[968] = 3'b0;
        for (loop_968 = 0; loop_968 < NUM_CELL; loop_968++) begin
         if ({b[8],a[30]}) == loop_968[1:0]) begin
          match_flag_968 = 1'b1;
          addr[968] = loop_968[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_969 = 1'b0;
        addr[969] = 3'b0;
        for (loop_969 = 0; loop_969 < NUM_CELL; loop_969++) begin
         if ({b[9],a[30]}) == loop_969[1:0]) begin
          match_flag_969 = 1'b1;
          addr[969] = loop_969[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_970 = 1'b0;
        addr[970] = 3'b0;
        for (loop_970 = 0; loop_970 < NUM_CELL; loop_970++) begin
         if ({b[10],a[30]}) == loop_970[1:0]) begin
          match_flag_970 = 1'b1;
          addr[970] = loop_970[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_971 = 1'b0;
        addr[971] = 3'b0;
        for (loop_971 = 0; loop_971 < NUM_CELL; loop_971++) begin
         if ({b[11],a[30]}) == loop_971[1:0]) begin
          match_flag_971 = 1'b1;
          addr[971] = loop_971[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_972 = 1'b0;
        addr[972] = 3'b0;
        for (loop_972 = 0; loop_972 < NUM_CELL; loop_972++) begin
         if ({b[12],a[30]}) == loop_972[1:0]) begin
          match_flag_972 = 1'b1;
          addr[972] = loop_972[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_973 = 1'b0;
        addr[973] = 3'b0;
        for (loop_973 = 0; loop_973 < NUM_CELL; loop_973++) begin
         if ({b[13],a[30]}) == loop_973[1:0]) begin
          match_flag_973 = 1'b1;
          addr[973] = loop_973[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_974 = 1'b0;
        addr[974] = 3'b0;
        for (loop_974 = 0; loop_974 < NUM_CELL; loop_974++) begin
         if ({b[14],a[30]}) == loop_974[1:0]) begin
          match_flag_974 = 1'b1;
          addr[974] = loop_974[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_975 = 1'b0;
        addr[975] = 3'b0;
        for (loop_975 = 0; loop_975 < NUM_CELL; loop_975++) begin
         if ({b[15],a[30]}) == loop_975[1:0]) begin
          match_flag_975 = 1'b1;
          addr[975] = loop_975[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_976 = 1'b0;
        addr[976] = 3'b0;
        for (loop_976 = 0; loop_976 < NUM_CELL; loop_976++) begin
         if ({b[16],a[30]}) == loop_976[1:0]) begin
          match_flag_976 = 1'b1;
          addr[976] = loop_976[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_977 = 1'b0;
        addr[977] = 3'b0;
        for (loop_977 = 0; loop_977 < NUM_CELL; loop_977++) begin
         if ({b[17],a[30]}) == loop_977[1:0]) begin
          match_flag_977 = 1'b1;
          addr[977] = loop_977[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_978 = 1'b0;
        addr[978] = 3'b0;
        for (loop_978 = 0; loop_978 < NUM_CELL; loop_978++) begin
         if ({b[18],a[30]}) == loop_978[1:0]) begin
          match_flag_978 = 1'b1;
          addr[978] = loop_978[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_979 = 1'b0;
        addr[979] = 3'b0;
        for (loop_979 = 0; loop_979 < NUM_CELL; loop_979++) begin
         if ({b[19],a[30]}) == loop_979[1:0]) begin
          match_flag_979 = 1'b1;
          addr[979] = loop_979[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_980 = 1'b0;
        addr[980] = 3'b0;
        for (loop_980 = 0; loop_980 < NUM_CELL; loop_980++) begin
         if ({b[20],a[30]}) == loop_980[1:0]) begin
          match_flag_980 = 1'b1;
          addr[980] = loop_980[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_981 = 1'b0;
        addr[981] = 3'b0;
        for (loop_981 = 0; loop_981 < NUM_CELL; loop_981++) begin
         if ({b[21],a[30]}) == loop_981[1:0]) begin
          match_flag_981 = 1'b1;
          addr[981] = loop_981[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_982 = 1'b0;
        addr[982] = 3'b0;
        for (loop_982 = 0; loop_982 < NUM_CELL; loop_982++) begin
         if ({b[22],a[30]}) == loop_982[1:0]) begin
          match_flag_982 = 1'b1;
          addr[982] = loop_982[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_983 = 1'b0;
        addr[983] = 3'b0;
        for (loop_983 = 0; loop_983 < NUM_CELL; loop_983++) begin
         if ({b[23],a[30]}) == loop_983[1:0]) begin
          match_flag_983 = 1'b1;
          addr[983] = loop_983[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_984 = 1'b0;
        addr[984] = 3'b0;
        for (loop_984 = 0; loop_984 < NUM_CELL; loop_984++) begin
         if ({b[24],a[30]}) == loop_984[1:0]) begin
          match_flag_984 = 1'b1;
          addr[984] = loop_984[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_985 = 1'b0;
        addr[985] = 3'b0;
        for (loop_985 = 0; loop_985 < NUM_CELL; loop_985++) begin
         if ({b[25],a[30]}) == loop_985[1:0]) begin
          match_flag_985 = 1'b1;
          addr[985] = loop_985[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_986 = 1'b0;
        addr[986] = 3'b0;
        for (loop_986 = 0; loop_986 < NUM_CELL; loop_986++) begin
         if ({b[26],a[30]}) == loop_986[1:0]) begin
          match_flag_986 = 1'b1;
          addr[986] = loop_986[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_987 = 1'b0;
        addr[987] = 3'b0;
        for (loop_987 = 0; loop_987 < NUM_CELL; loop_987++) begin
         if ({b[27],a[30]}) == loop_987[1:0]) begin
          match_flag_987 = 1'b1;
          addr[987] = loop_987[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_988 = 1'b0;
        addr[988] = 3'b0;
        for (loop_988 = 0; loop_988 < NUM_CELL; loop_988++) begin
         if ({b[28],a[30]}) == loop_988[1:0]) begin
          match_flag_988 = 1'b1;
          addr[988] = loop_988[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_989 = 1'b0;
        addr[989] = 3'b0;
        for (loop_989 = 0; loop_989 < NUM_CELL; loop_989++) begin
         if ({b[29],a[30]}) == loop_989[1:0]) begin
          match_flag_989 = 1'b1;
          addr[989] = loop_989[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_990 = 1'b0;
        addr[990] = 3'b0;
        for (loop_990 = 0; loop_990 < NUM_CELL; loop_990++) begin
         if ({b[30],a[30]}) == loop_990[1:0]) begin
          match_flag_990 = 1'b1;
          addr[990] = loop_990[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_991 = 1'b0;
        addr[991] = 3'b0;
        for (loop_991 = 0; loop_991 < NUM_CELL; loop_991++) begin
         if ({b[31],a[30]}) == loop_991[1:0]) begin
          match_flag_991 = 1'b1;
          addr[991] = loop_991[1:0];
          break;
        end
      end
    end
    
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_992 = 1'b0;
        addr[992] = 3'b0;
        for (loop_992 = 0; loop_992 < NUM_CELL; loop_992++) begin
         if ({b[0],a[31]}) == loop_992[1:0]) begin
          match_flag_992 = 1'b1;
          addr[992] = loop_992[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_993 = 1'b0;
        addr[993] = 3'b0;
        for (loop_993 = 0; loop_993 < NUM_CELL; loop_993++) begin
         if ({b[1],a[31]}) == loop_993[1:0]) begin
          match_flag_993 = 1'b1;
          addr[993] = loop_993[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_994 = 1'b0;
        addr[994] = 3'b0;
        for (loop_994 = 0; loop_994 < NUM_CELL; loop_994++) begin
         if ({b[2],a[31]}) == loop_994[1:0]) begin
          match_flag_994 = 1'b1;
          addr[994] = loop_994[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_995 = 1'b0;
        addr[995] = 3'b0;
        for (loop_995 = 0; loop_995 < NUM_CELL; loop_995++) begin
         if ({b[3],a[31]}) == loop_995[1:0]) begin
          match_flag_995 = 1'b1;
          addr[995] = loop_995[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_996 = 1'b0;
        addr[996] = 3'b0;
        for (loop_996 = 0; loop_996 < NUM_CELL; loop_996++) begin
         if ({b[4],a[31]}) == loop_996[1:0]) begin
          match_flag_996 = 1'b1;
          addr[996] = loop_996[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_997 = 1'b0;
        addr[997] = 3'b0;
        for (loop_997 = 0; loop_997 < NUM_CELL; loop_997++) begin
         if ({b[5],a[31]}) == loop_997[1:0]) begin
          match_flag_997 = 1'b1;
          addr[997] = loop_997[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_998 = 1'b0;
        addr[998] = 3'b0;
        for (loop_998 = 0; loop_998 < NUM_CELL; loop_998++) begin
         if ({b[6],a[31]}) == loop_998[1:0]) begin
          match_flag_998 = 1'b1;
          addr[998] = loop_998[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_999 = 1'b0;
        addr[999] = 3'b0;
        for (loop_999 = 0; loop_999 < NUM_CELL; loop_999++) begin
         if ({b[7],a[31]}) == loop_999[1:0]) begin
          match_flag_999 = 1'b1;
          addr[999] = loop_999[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1000 = 1'b0;
        addr[1000] = 3'b0;
        for (loop_1000 = 0; loop_1000 < NUM_CELL; loop_1000++) begin
         if ({b[8],a[31]}) == loop_1000[1:0]) begin
          match_flag_1000 = 1'b1;
          addr[1000] = loop_1000[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1001 = 1'b0;
        addr[1001] = 3'b0;
        for (loop_1001 = 0; loop_1001 < NUM_CELL; loop_1001++) begin
         if ({b[9],a[31]}) == loop_1001[1:0]) begin
          match_flag_1001 = 1'b1;
          addr[1001] = loop_1001[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1002 = 1'b0;
        addr[1002] = 3'b0;
        for (loop_1002 = 0; loop_1002 < NUM_CELL; loop_1002++) begin
         if ({b[10],a[31]}) == loop_1002[1:0]) begin
          match_flag_1002 = 1'b1;
          addr[1002] = loop_1002[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1003 = 1'b0;
        addr[1003] = 3'b0;
        for (loop_1003 = 0; loop_1003 < NUM_CELL; loop_1003++) begin
         if ({b[11],a[31]}) == loop_1003[1:0]) begin
          match_flag_1003 = 1'b1;
          addr[1003] = loop_1003[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1004 = 1'b0;
        addr[1004] = 3'b0;
        for (loop_1004 = 0; loop_1004 < NUM_CELL; loop_1004++) begin
         if ({b[12],a[31]}) == loop_1004[1:0]) begin
          match_flag_1004 = 1'b1;
          addr[1004] = loop_1004[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1005 = 1'b0;
        addr[1005] = 3'b0;
        for (loop_1005 = 0; loop_1005 < NUM_CELL; loop_1005++) begin
         if ({b[13],a[31]}) == loop_1005[1:0]) begin
          match_flag_1005 = 1'b1;
          addr[1005] = loop_1005[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1006 = 1'b0;
        addr[1006] = 3'b0;
        for (loop_1006 = 0; loop_1006 < NUM_CELL; loop_1006++) begin
         if ({b[14],a[31]}) == loop_1006[1:0]) begin
          match_flag_1006 = 1'b1;
          addr[1006] = loop_1006[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1007 = 1'b0;
        addr[1007] = 3'b0;
        for (loop_1007 = 0; loop_1007 < NUM_CELL; loop_1007++) begin
         if ({b[15],a[31]}) == loop_1007[1:0]) begin
          match_flag_1007 = 1'b1;
          addr[1007] = loop_1007[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1008 = 1'b0;
        addr[1008] = 3'b0;
        for (loop_1008 = 0; loop_1008 < NUM_CELL; loop_1008++) begin
         if ({b[16],a[31]}) == loop_1008[1:0]) begin
          match_flag_1008 = 1'b1;
          addr[1008] = loop_1008[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1009 = 1'b0;
        addr[1009] = 3'b0;
        for (loop_1009 = 0; loop_1009 < NUM_CELL; loop_1009++) begin
         if ({b[17],a[31]}) == loop_1009[1:0]) begin
          match_flag_1009 = 1'b1;
          addr[1009] = loop_1009[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1010 = 1'b0;
        addr[1010] = 3'b0;
        for (loop_1010 = 0; loop_1010 < NUM_CELL; loop_1010++) begin
         if ({b[18],a[31]}) == loop_1010[1:0]) begin
          match_flag_1010 = 1'b1;
          addr[1010] = loop_1010[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1011 = 1'b0;
        addr[1011] = 3'b0;
        for (loop_1011 = 0; loop_1011 < NUM_CELL; loop_1011++) begin
         if ({b[19],a[31]}) == loop_1011[1:0]) begin
          match_flag_1011 = 1'b1;
          addr[1011] = loop_1011[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1012 = 1'b0;
        addr[1012] = 3'b0;
        for (loop_1012 = 0; loop_1012 < NUM_CELL; loop_1012++) begin
         if ({b[20],a[31]}) == loop_1012[1:0]) begin
          match_flag_1012 = 1'b1;
          addr[1012] = loop_1012[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1013 = 1'b0;
        addr[1013] = 3'b0;
        for (loop_1013 = 0; loop_1013 < NUM_CELL; loop_1013++) begin
         if ({b[21],a[31]}) == loop_1013[1:0]) begin
          match_flag_1013 = 1'b1;
          addr[1013] = loop_1013[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1014 = 1'b0;
        addr[1014] = 3'b0;
        for (loop_1014 = 0; loop_1014 < NUM_CELL; loop_1014++) begin
         if ({b[22],a[31]}) == loop_1014[1:0]) begin
          match_flag_1014 = 1'b1;
          addr[1014] = loop_1014[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1015 = 1'b0;
        addr[1015] = 3'b0;
        for (loop_1015 = 0; loop_1015 < NUM_CELL; loop_1015++) begin
         if ({b[23],a[31]}) == loop_1015[1:0]) begin
          match_flag_1015 = 1'b1;
          addr[1015] = loop_1015[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1016 = 1'b0;
        addr[1016] = 3'b0;
        for (loop_1016 = 0; loop_1016 < NUM_CELL; loop_1016++) begin
         if ({b[24],a[31]}) == loop_1016[1:0]) begin
          match_flag_1016 = 1'b1;
          addr[1016] = loop_1016[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1017 = 1'b0;
        addr[1017] = 3'b0;
        for (loop_1017 = 0; loop_1017 < NUM_CELL; loop_1017++) begin
         if ({b[25],a[31]}) == loop_1017[1:0]) begin
          match_flag_1017 = 1'b1;
          addr[1017] = loop_1017[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1018 = 1'b0;
        addr[1018] = 3'b0;
        for (loop_1018 = 0; loop_1018 < NUM_CELL; loop_1018++) begin
         if ({b[26],a[31]}) == loop_1018[1:0]) begin
          match_flag_1018 = 1'b1;
          addr[1018] = loop_1018[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1019 = 1'b0;
        addr[1019] = 3'b0;
        for (loop_1019 = 0; loop_1019 < NUM_CELL; loop_1019++) begin
         if ({b[27],a[31]}) == loop_1019[1:0]) begin
          match_flag_1019 = 1'b1;
          addr[1019] = loop_1019[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1020 = 1'b0;
        addr[1020] = 3'b0;
        for (loop_1020 = 0; loop_1020 < NUM_CELL; loop_1020++) begin
         if ({b[28],a[31]}) == loop_1020[1:0]) begin
          match_flag_1020 = 1'b1;
          addr[1020] = loop_1020[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1021 = 1'b0;
        addr[1021] = 3'b0;
        for (loop_1021 = 0; loop_1021 < NUM_CELL; loop_1021++) begin
         if ({b[29],a[31]}) == loop_1021[1:0]) begin
          match_flag_1021 = 1'b1;
          addr[1021] = loop_1021[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1022 = 1'b0;
        addr[1022] = 3'b0;
        for (loop_1022 = 0; loop_1022 < NUM_CELL; loop_1022++) begin
         if ({b[30],a[31]}) == loop_1022[1:0]) begin
          match_flag_1022 = 1'b1;
          addr[1022] = loop_1022[1:0];
          break;
        end
      end
    end
     always_ff @(posedge clk) begin
      if (data_flag) begin
        match_flag_1023 = 1'b0;
        addr[1023] = 3'b0;
        for (loop_1023 = 0; loop_1023 < NUM_CELL; loop_1023++) begin
         if ({b[31],a[31]}) == loop_1023[1:0]) begin
          match_flag_1023 = 1'b1;
          addr[1023] = loop_1023[1:0];
          break;
        end
      end
    end

 
endmodule
